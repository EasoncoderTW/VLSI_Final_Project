module chip(
//inputs
    PI_clk,
    PI_rst,
    PI_Inst_Cahe_readAddr_ready,
    PI_Inst_Cahe_readData_data,
    PI_Inst_Cahe_readData_valid,
    PI_Inst_Cahe_writeAddr_ready,
    PI_Inst_Cahe_writeData_ready,
    PI_Inst_Cahe_writeResp_msg,
    PI_Inst_Cahe_writeResp_valid,
    PI_Data_Cahe_readAddr_ready,
    PI_Data_Cahe_readData_data,
    PI_Data_Cahe_readData_valid,
    PI_Data_Cahe_writeAddr_ready,
    PI_Data_Cahe_writeData_ready,
    PI_Data_Cahe_writeResp_msg,
    PI_Data_Cahe_writeResp_valid,
//outputs
    PO_Inst_Cahe_readAddr_addr,
    PO_Inst_Cahe_readAddr_valid,
    PO_Inst_Cahe_readData_ready,
    PO_Inst_Cahe_writeAddr_addr,
    PO_Inst_Cahe_writeAddr_valid,
    PO_Inst_Cahe_writeData_data,
    PO_Inst_Cahe_writeData_strb,
    PO_Inst_Cahe_writeData_valid,
    PO_Inst_Cahe_writeResp_ready,
    PO_Data_Cahe_readAddr_addr,
    PO_Data_Cahe_readAddr_valid,
    PO_Data_Cahe_readData_ready,
    PO_Data_Cahe_writeAddr_addr,
    PO_Data_Cahe_writeAddr_valid,
    PO_Data_Cahe_writeData_data,
    PO_Data_Cahe_writeData_strb,
    PO_Data_Cahe_writeData_valid,
    PO_Data_Cahe_writeResp_ready,
    PO_halt
);
    input            PI_clk;                       //0
    input            PI_rst;                       //0
    input            PI_Inst_Cahe_readAddr_ready;  //0
    input   [127:0]  PI_Inst_Cahe_readData_data;   //0
    input            PI_Inst_Cahe_readData_valid;  //0
    input            PI_Inst_Cahe_writeAddr_ready; //0
    input            PI_Inst_Cahe_writeData_ready; //0
    input   [31:0]   PI_Inst_Cahe_writeResp_msg;   //0
    input            PI_Inst_Cahe_writeResp_valid; //0
    input            PI_Data_Cahe_readAddr_ready;  //2
    input   [127:0]  PI_Data_Cahe_readData_data;   //2
    input            PI_Data_Cahe_readData_valid;  //2
    input            PI_Data_Cahe_writeAddr_ready; //2
    input            PI_Data_Cahe_writeData_ready; //2
    input   [31:0]   PI_Data_Cahe_writeResp_msg;   //2
    input            PI_Data_Cahe_writeResp_valid; //2
    
    output  [31:0]   PO_Inst_Cahe_readAddr_addr;   //1
    output           PO_Inst_Cahe_readAddr_valid;  //1
    output           PO_Inst_Cahe_readData_ready;  //1
    output  [31:0]   PO_Inst_Cahe_writeAddr_addr;  //1
    output           PO_Inst_Cahe_writeAddr_valid; //1
    output  [127:0]  PO_Inst_Cahe_writeData_data;  //1 
    output  [15:0]   PO_Inst_Cahe_writeData_strb;  //1
    output           PO_Inst_Cahe_writeData_valid; //1
    output           PO_Inst_Cahe_writeResp_ready; //1
    output  [31:0]   PO_Data_Cahe_readAddr_addr;   //3
    output           PO_Data_Cahe_readAddr_valid;  //3
    output           PO_Data_Cahe_readData_ready;  //3
    output  [31:0]   PO_Data_Cahe_writeAddr_addr;  //3
    output           PO_Data_Cahe_writeAddr_valid; //3
    output  [127:0]  PO_Data_Cahe_writeData_data;  //3  
    output  [15:0]   PO_Data_Cahe_writeData_strb;  //3
    output           PO_Data_Cahe_writeData_valid; //3
    output           PO_Data_Cahe_writeResp_ready; //3
    output           PO_halt;                      //0

    wire             WIRE_clk;
    wire             WIRE_rst;
    wire             WIRE_Inst_Cahe_readAddr_ready;
    wire   [127:0]   WIRE_Inst_Cahe_readData_data;
    wire             WIRE_Inst_Cahe_readData_valid;
    wire             WIRE_Inst_Cahe_writeAddr_ready;
    wire             WIRE_Inst_Cahe_writeData_ready;
    wire   [31:0]    WIRE_Inst_Cahe_writeResp_msg;
    wire             WIRE_Inst_Cahe_writeResp_valid;
    wire             WIRE_Data_Cahe_readAddr_ready;
    wire   [127:0]   WIRE_Data_Cahe_readData_data;
    wire             WIRE_Data_Cahe_readData_valid;
    wire             WIRE_Data_Cahe_writeAddr_ready;
    wire             WIRE_Data_Cahe_writeData_ready;
    wire   [31:0]    WIRE_Data_Cahe_writeResp_msg;
    wire             WIRE_Data_Cahe_writeResp_valid;
    wire  [31:0]     WIRE_Inst_Cahe_readAddr_addr;
    wire             WIRE_Inst_Cahe_readAddr_valid;
    wire             WIRE_Inst_Cahe_readData_ready;
    wire  [31:0]     WIRE_Inst_Cahe_writeAddr_addr;
    wire             WIRE_Inst_Cahe_writeAddr_valid;
    wire  [127:0]    WIRE_Inst_Cahe_writeData_data;
    wire  [15:0]     WIRE_Inst_Cahe_writeData_strb;
    wire             WIRE_Inst_Cahe_writeData_valid;
    wire             WIRE_Inst_Cahe_writeResp_ready;
    wire  [31:0]     WIRE_Data_Cahe_readAddr_addr;
    wire             WIRE_Data_Cahe_readAddr_valid;
    wire             WIRE_Data_Cahe_readData_ready;
    wire  [31:0]     WIRE_Data_Cahe_writeAddr_addr;
    wire             WIRE_Data_Cahe_writeAddr_valid;
    wire  [127:0]    WIRE_Data_Cahe_writeData_data;
    wire  [15:0]     WIRE_Data_Cahe_writeData_strb;
    wire             WIRE_Data_Cahe_writeData_valid;
    wire             WIRE_Data_Cahe_writeResp_ready;
    wire             WIRE_halt;

CPU CPU(
    .clk(WIRE_clk)
    .rst(WIRE_rst)
    .Inst_Cahe_readAddr_ready(WIRE_Inst_Cahe_readAddr_ready)
    .Inst_Cahe_readData_data(WIRE_Inst_Cahe_readData_data)
    .Inst_Cahe_readData_valid(WIRE_Inst_Cahe_readData_valid)
    .Inst_Cahe_writeAddr_ready(WIRE_Inst_Cahe_writeAddr_ready)
    .Inst_Cahe_writeData_ready(WIRE_Inst_Cahe_writeData_ready)
    .Inst_Cahe_writeResp_msg(WIRE_Inst_Cahe_writeResp_msg)
    .Inst_Cahe_writeResp_valid(WIRE_Inst_Cahe_writeResp_valid)
    .Data_Cahe_readAddr_ready(WIRE_Data_Cahe_readAddr_ready)
    .Data_Cahe_readData_data(WIRE_Data_Cahe_readData_data)
    .Data_Cahe_readData_valid(WIRE_Data_Cahe_readData_valid)
    .Data_Cahe_writeAddr_ready(WIRE_Data_Cahe_writeAddr_ready)
    .Data_Cahe_writeData_ready(WIRE_Data_Cahe_writeData_ready)
    .Data_Cahe_writeResp_msg(WIRE_Data_Cahe_writeResp_msg)
    .Data_Cahe_writeResp_valid(WIRE_Data_Cahe_writeResp_valid)
    .Inst_Cahe_readAddr_addr(WIRE_Inst_Cahe_readAddr_addr)
    .Inst_Cahe_readAddr_valid(WIRE_Inst_Cahe_readAddr_valid)
    .Inst_Cahe_readData_ready(WIRE_Inst_Cahe_readData_ready)
    .Inst_Cahe_writeAddr_addr(WIRE_Inst_Cahe_writeAddr_addr)
    .Inst_Cahe_writeAddr_valid(WIRE_Inst_Cahe_writeAddr_valid)
    .Inst_Cahe_writeData_data(WIRE_Inst_Cahe_writeData_data)
    .Inst_Cahe_writeData_strb(WIRE_Inst_Cahe_writeData_strb)
    .Inst_Cahe_writeData_valid(WIRE_Inst_Cahe_writeData_valid)
    .Inst_Cahe_writeResp_ready(WIRE_Inst_Cahe_writeResp_ready)
    .Data_Cahe_readAddr_addr(WIRE_Data_Cahe_readAddr_addr)
    .Data_Cahe_readAddr_valid(WIRE_Data_Cahe_readAddr_valid)
    .Data_Cahe_readData_ready(WIRE_Data_Cahe_readData_ready)
    .Data_Cahe_writeAddr_addr(WIRE_Data_Cahe_writeAddr_addr)
    .Data_Cahe_writeAddr_valid(WIRE_Data_Cahe_writeAddr_valid)
    .Data_Cahe_writeData_data(WIRE_Data_Cahe_writeData_data)
    .Data_Cahe_writeData_strb(WIRE_Data_Cahe_writeData_strb)
    .Data_Cahe_writeData_valid(WIRE_Data_Cahe_writeData_valid)
    .Data_Cahe_writeResp_ready(WIRE_Data_Cahe_writeResp_ready)
    .halt(WIRE_halt)
);

// input pads: PDIDGZ (.PAD(PI), .C(WIRE))
// CORNER0
PDIDGZ PAD_Inst_Cahe_readAddr_ready   (.PAD(PI_Inst_Cahe_readAddr_ready), .C(WIRE_Inst_Cahe_readAddr_ready));

PDIDGZ PAD_Inst_Cahe_readData_data0 (.PAD(PI_Inst_Cahe_readData_data[0]), .C(WIRE_Inst_Cahe_readData_data[0]));
PDIDGZ PAD_Inst_Cahe_readData_data1 (.PAD(PI_Inst_Cahe_readData_data[1]), .C(WIRE_Inst_Cahe_readData_data[1]));
PDIDGZ PAD_Inst_Cahe_readData_data2 (.PAD(PI_Inst_Cahe_readData_data[2]), .C(WIRE_Inst_Cahe_readData_data[2]));
PDIDGZ PAD_Inst_Cahe_readData_data3 (.PAD(PI_Inst_Cahe_readData_data[3]), .C(WIRE_Inst_Cahe_readData_data[3]));
PDIDGZ PAD_Inst_Cahe_readData_data4 (.PAD(PI_Inst_Cahe_readData_data[4]), .C(WIRE_Inst_Cahe_readData_data[4]));
PDIDGZ PAD_Inst_Cahe_readData_data5 (.PAD(PI_Inst_Cahe_readData_data[5]), .C(WIRE_Inst_Cahe_readData_data[5]));
PDIDGZ PAD_Inst_Cahe_readData_data6 (.PAD(PI_Inst_Cahe_readData_data[6]), .C(WIRE_Inst_Cahe_readData_data[6]));
PDIDGZ PAD_Inst_Cahe_readData_data7 (.PAD(PI_Inst_Cahe_readData_data[7]), .C(WIRE_Inst_Cahe_readData_data[7]));
PDIDGZ PAD_Inst_Cahe_readData_data8 (.PAD(PI_Inst_Cahe_readData_data[8]), .C(WIRE_Inst_Cahe_readData_data[8]));
PDIDGZ PAD_Inst_Cahe_readData_data9 (.PAD(PI_Inst_Cahe_readData_data[9]), .C(WIRE_Inst_Cahe_readData_data[9]));
PDIDGZ PAD_Inst_Cahe_readData_data10 (.PAD(PI_Inst_Cahe_readData_data[10]), .C(WIRE_Inst_Cahe_readData_data[10]));
PDIDGZ PAD_Inst_Cahe_readData_data11 (.PAD(PI_Inst_Cahe_readData_data[11]), .C(WIRE_Inst_Cahe_readData_data[11]));
PDIDGZ PAD_Inst_Cahe_readData_data12 (.PAD(PI_Inst_Cahe_readData_data[12]), .C(WIRE_Inst_Cahe_readData_data[12]));
PDIDGZ PAD_Inst_Cahe_readData_data13 (.PAD(PI_Inst_Cahe_readData_data[13]), .C(WIRE_Inst_Cahe_readData_data[13]));
PDIDGZ PAD_Inst_Cahe_readData_data14 (.PAD(PI_Inst_Cahe_readData_data[14]), .C(WIRE_Inst_Cahe_readData_data[14]));
PDIDGZ PAD_Inst_Cahe_readData_data15 (.PAD(PI_Inst_Cahe_readData_data[15]), .C(WIRE_Inst_Cahe_readData_data[15]));
PDIDGZ PAD_Inst_Cahe_readData_data16 (.PAD(PI_Inst_Cahe_readData_data[16]), .C(WIRE_Inst_Cahe_readData_data[16]));
PDIDGZ PAD_Inst_Cahe_readData_data17 (.PAD(PI_Inst_Cahe_readData_data[17]), .C(WIRE_Inst_Cahe_readData_data[17]));
PDIDGZ PAD_Inst_Cahe_readData_data18 (.PAD(PI_Inst_Cahe_readData_data[18]), .C(WIRE_Inst_Cahe_readData_data[18]));
PDIDGZ PAD_Inst_Cahe_readData_data19 (.PAD(PI_Inst_Cahe_readData_data[19]), .C(WIRE_Inst_Cahe_readData_data[19]));
PDIDGZ PAD_Inst_Cahe_readData_data20 (.PAD(PI_Inst_Cahe_readData_data[20]), .C(WIRE_Inst_Cahe_readData_data[20]));
PDIDGZ PAD_Inst_Cahe_readData_data21 (.PAD(PI_Inst_Cahe_readData_data[21]), .C(WIRE_Inst_Cahe_readData_data[21]));
PDIDGZ PAD_Inst_Cahe_readData_data22 (.PAD(PI_Inst_Cahe_readData_data[22]), .C(WIRE_Inst_Cahe_readData_data[22]));
PDIDGZ PAD_Inst_Cahe_readData_data23 (.PAD(PI_Inst_Cahe_readData_data[23]), .C(WIRE_Inst_Cahe_readData_data[23]));
PDIDGZ PAD_Inst_Cahe_readData_data24 (.PAD(PI_Inst_Cahe_readData_data[24]), .C(WIRE_Inst_Cahe_readData_data[24]));
PDIDGZ PAD_Inst_Cahe_readData_data25 (.PAD(PI_Inst_Cahe_readData_data[25]), .C(WIRE_Inst_Cahe_readData_data[25]));
PDIDGZ PAD_Inst_Cahe_readData_data26 (.PAD(PI_Inst_Cahe_readData_data[26]), .C(WIRE_Inst_Cahe_readData_data[26]));
PDIDGZ PAD_Inst_Cahe_readData_data27 (.PAD(PI_Inst_Cahe_readData_data[27]), .C(WIRE_Inst_Cahe_readData_data[27]));
PDIDGZ PAD_Inst_Cahe_readData_data28 (.PAD(PI_Inst_Cahe_readData_data[28]), .C(WIRE_Inst_Cahe_readData_data[28]));
PDIDGZ PAD_Inst_Cahe_readData_data29 (.PAD(PI_Inst_Cahe_readData_data[29]), .C(WIRE_Inst_Cahe_readData_data[29]));
PDIDGZ PAD_Inst_Cahe_readData_data30 (.PAD(PI_Inst_Cahe_readData_data[30]), .C(WIRE_Inst_Cahe_readData_data[30]));
PDIDGZ PAD_Inst_Cahe_readData_data31 (.PAD(PI_Inst_Cahe_readData_data[31]), .C(WIRE_Inst_Cahe_readData_data[31]));
PDIDGZ PAD_Inst_Cahe_readData_data32 (.PAD(PI_Inst_Cahe_readData_data[32]), .C(WIRE_Inst_Cahe_readData_data[32]));
PDIDGZ PAD_Inst_Cahe_readData_data33 (.PAD(PI_Inst_Cahe_readData_data[33]), .C(WIRE_Inst_Cahe_readData_data[33]));
PDIDGZ PAD_Inst_Cahe_readData_data34 (.PAD(PI_Inst_Cahe_readData_data[34]), .C(WIRE_Inst_Cahe_readData_data[34]));
PDIDGZ PAD_Inst_Cahe_readData_data35 (.PAD(PI_Inst_Cahe_readData_data[35]), .C(WIRE_Inst_Cahe_readData_data[35]));
PDIDGZ PAD_Inst_Cahe_readData_data36 (.PAD(PI_Inst_Cahe_readData_data[36]), .C(WIRE_Inst_Cahe_readData_data[36]));
PDIDGZ PAD_Inst_Cahe_readData_data37 (.PAD(PI_Inst_Cahe_readData_data[37]), .C(WIRE_Inst_Cahe_readData_data[37]));
PDIDGZ PAD_Inst_Cahe_readData_data38 (.PAD(PI_Inst_Cahe_readData_data[38]), .C(WIRE_Inst_Cahe_readData_data[38]));
PDIDGZ PAD_Inst_Cahe_readData_data39 (.PAD(PI_Inst_Cahe_readData_data[39]), .C(WIRE_Inst_Cahe_readData_data[39]));
PDIDGZ PAD_Inst_Cahe_readData_data40 (.PAD(PI_Inst_Cahe_readData_data[40]), .C(WIRE_Inst_Cahe_readData_data[40]));
PDIDGZ PAD_Inst_Cahe_readData_data41 (.PAD(PI_Inst_Cahe_readData_data[41]), .C(WIRE_Inst_Cahe_readData_data[41]));
PDIDGZ PAD_Inst_Cahe_readData_data42 (.PAD(PI_Inst_Cahe_readData_data[42]), .C(WIRE_Inst_Cahe_readData_data[42]));
PDIDGZ PAD_Inst_Cahe_readData_data43 (.PAD(PI_Inst_Cahe_readData_data[43]), .C(WIRE_Inst_Cahe_readData_data[43]));
PDIDGZ PAD_Inst_Cahe_readData_data44 (.PAD(PI_Inst_Cahe_readData_data[44]), .C(WIRE_Inst_Cahe_readData_data[44]));
PDIDGZ PAD_Inst_Cahe_readData_data45 (.PAD(PI_Inst_Cahe_readData_data[45]), .C(WIRE_Inst_Cahe_readData_data[45]));
PDIDGZ PAD_Inst_Cahe_readData_data46 (.PAD(PI_Inst_Cahe_readData_data[46]), .C(WIRE_Inst_Cahe_readData_data[46]));
PDIDGZ PAD_Inst_Cahe_readData_data47 (.PAD(PI_Inst_Cahe_readData_data[47]), .C(WIRE_Inst_Cahe_readData_data[47]));
PDIDGZ PAD_Inst_Cahe_readData_data48 (.PAD(PI_Inst_Cahe_readData_data[48]), .C(WIRE_Inst_Cahe_readData_data[48]));
PDIDGZ PAD_Inst_Cahe_readData_data49 (.PAD(PI_Inst_Cahe_readData_data[49]), .C(WIRE_Inst_Cahe_readData_data[49]));
PDIDGZ PAD_Inst_Cahe_readData_data50 (.PAD(PI_Inst_Cahe_readData_data[50]), .C(WIRE_Inst_Cahe_readData_data[50]));
PDIDGZ PAD_Inst_Cahe_readData_data51 (.PAD(PI_Inst_Cahe_readData_data[51]), .C(WIRE_Inst_Cahe_readData_data[51]));
PDIDGZ PAD_Inst_Cahe_readData_data52 (.PAD(PI_Inst_Cahe_readData_data[52]), .C(WIRE_Inst_Cahe_readData_data[52]));
PDIDGZ PAD_Inst_Cahe_readData_data53 (.PAD(PI_Inst_Cahe_readData_data[53]), .C(WIRE_Inst_Cahe_readData_data[53]));
PDIDGZ PAD_Inst_Cahe_readData_data54 (.PAD(PI_Inst_Cahe_readData_data[54]), .C(WIRE_Inst_Cahe_readData_data[54]));
PDIDGZ PAD_Inst_Cahe_readData_data55 (.PAD(PI_Inst_Cahe_readData_data[55]), .C(WIRE_Inst_Cahe_readData_data[55]));
PDIDGZ PAD_Inst_Cahe_readData_data56 (.PAD(PI_Inst_Cahe_readData_data[56]), .C(WIRE_Inst_Cahe_readData_data[56]));
PDIDGZ PAD_Inst_Cahe_readData_data57 (.PAD(PI_Inst_Cahe_readData_data[57]), .C(WIRE_Inst_Cahe_readData_data[57]));
PDIDGZ PAD_Inst_Cahe_readData_data58 (.PAD(PI_Inst_Cahe_readData_data[58]), .C(WIRE_Inst_Cahe_readData_data[58]));
PDIDGZ PAD_Inst_Cahe_readData_data59 (.PAD(PI_Inst_Cahe_readData_data[59]), .C(WIRE_Inst_Cahe_readData_data[59]));
PDIDGZ PAD_Inst_Cahe_readData_data60 (.PAD(PI_Inst_Cahe_readData_data[60]), .C(WIRE_Inst_Cahe_readData_data[60]));
PDIDGZ PAD_Inst_Cahe_readData_data61 (.PAD(PI_Inst_Cahe_readData_data[61]), .C(WIRE_Inst_Cahe_readData_data[61]));
PDIDGZ PAD_Inst_Cahe_readData_data62 (.PAD(PI_Inst_Cahe_readData_data[62]), .C(WIRE_Inst_Cahe_readData_data[62]));
PDIDGZ PAD_Inst_Cahe_readData_data63 (.PAD(PI_Inst_Cahe_readData_data[63]), .C(WIRE_Inst_Cahe_readData_data[63]));
PDIDGZ PAD_Inst_Cahe_readData_data64 (.PAD(PI_Inst_Cahe_readData_data[64]), .C(WIRE_Inst_Cahe_readData_data[64]));
PDIDGZ PAD_Inst_Cahe_readData_data65 (.PAD(PI_Inst_Cahe_readData_data[65]), .C(WIRE_Inst_Cahe_readData_data[65]));
PDIDGZ PAD_Inst_Cahe_readData_data66 (.PAD(PI_Inst_Cahe_readData_data[66]), .C(WIRE_Inst_Cahe_readData_data[66]));
PDIDGZ PAD_Inst_Cahe_readData_data67 (.PAD(PI_Inst_Cahe_readData_data[67]), .C(WIRE_Inst_Cahe_readData_data[67]));
PDIDGZ PAD_Inst_Cahe_readData_data68 (.PAD(PI_Inst_Cahe_readData_data[68]), .C(WIRE_Inst_Cahe_readData_data[68]));
PDIDGZ PAD_Inst_Cahe_readData_data69 (.PAD(PI_Inst_Cahe_readData_data[69]), .C(WIRE_Inst_Cahe_readData_data[69]));
PDIDGZ PAD_Inst_Cahe_readData_data70 (.PAD(PI_Inst_Cahe_readData_data[70]), .C(WIRE_Inst_Cahe_readData_data[70]));
PDIDGZ PAD_Inst_Cahe_readData_data71 (.PAD(PI_Inst_Cahe_readData_data[71]), .C(WIRE_Inst_Cahe_readData_data[71]));
PDIDGZ PAD_Inst_Cahe_readData_data72 (.PAD(PI_Inst_Cahe_readData_data[72]), .C(WIRE_Inst_Cahe_readData_data[72]));
PDIDGZ PAD_Inst_Cahe_readData_data73 (.PAD(PI_Inst_Cahe_readData_data[73]), .C(WIRE_Inst_Cahe_readData_data[73]));
PDIDGZ PAD_Inst_Cahe_readData_data74 (.PAD(PI_Inst_Cahe_readData_data[74]), .C(WIRE_Inst_Cahe_readData_data[74]));
PDIDGZ PAD_Inst_Cahe_readData_data75 (.PAD(PI_Inst_Cahe_readData_data[75]), .C(WIRE_Inst_Cahe_readData_data[75]));
PDIDGZ PAD_Inst_Cahe_readData_data76 (.PAD(PI_Inst_Cahe_readData_data[76]), .C(WIRE_Inst_Cahe_readData_data[76]));
PDIDGZ PAD_Inst_Cahe_readData_data77 (.PAD(PI_Inst_Cahe_readData_data[77]), .C(WIRE_Inst_Cahe_readData_data[77]));
PDIDGZ PAD_Inst_Cahe_readData_data78 (.PAD(PI_Inst_Cahe_readData_data[78]), .C(WIRE_Inst_Cahe_readData_data[78]));
PDIDGZ PAD_Inst_Cahe_readData_data79 (.PAD(PI_Inst_Cahe_readData_data[79]), .C(WIRE_Inst_Cahe_readData_data[79]));
PDIDGZ PAD_Inst_Cahe_readData_data80 (.PAD(PI_Inst_Cahe_readData_data[80]), .C(WIRE_Inst_Cahe_readData_data[80]));
PDIDGZ PAD_Inst_Cahe_readData_data81 (.PAD(PI_Inst_Cahe_readData_data[81]), .C(WIRE_Inst_Cahe_readData_data[81]));
PDIDGZ PAD_Inst_Cahe_readData_data82 (.PAD(PI_Inst_Cahe_readData_data[82]), .C(WIRE_Inst_Cahe_readData_data[82]));
PDIDGZ PAD_Inst_Cahe_readData_data83 (.PAD(PI_Inst_Cahe_readData_data[83]), .C(WIRE_Inst_Cahe_readData_data[83]));
PDIDGZ PAD_Inst_Cahe_readData_data84 (.PAD(PI_Inst_Cahe_readData_data[84]), .C(WIRE_Inst_Cahe_readData_data[84]));
PDIDGZ PAD_Inst_Cahe_readData_data85 (.PAD(PI_Inst_Cahe_readData_data[85]), .C(WIRE_Inst_Cahe_readData_data[85]));
PDIDGZ PAD_Inst_Cahe_readData_data86 (.PAD(PI_Inst_Cahe_readData_data[86]), .C(WIRE_Inst_Cahe_readData_data[86]));
PDIDGZ PAD_Inst_Cahe_readData_data87 (.PAD(PI_Inst_Cahe_readData_data[87]), .C(WIRE_Inst_Cahe_readData_data[87]));
PDIDGZ PAD_Inst_Cahe_readData_data88 (.PAD(PI_Inst_Cahe_readData_data[88]), .C(WIRE_Inst_Cahe_readData_data[88]));
PDIDGZ PAD_Inst_Cahe_readData_data89 (.PAD(PI_Inst_Cahe_readData_data[89]), .C(WIRE_Inst_Cahe_readData_data[89]));
PDIDGZ PAD_Inst_Cahe_readData_data90 (.PAD(PI_Inst_Cahe_readData_data[90]), .C(WIRE_Inst_Cahe_readData_data[90]));
PDIDGZ PAD_Inst_Cahe_readData_data91 (.PAD(PI_Inst_Cahe_readData_data[91]), .C(WIRE_Inst_Cahe_readData_data[91]));
PDIDGZ PAD_Inst_Cahe_readData_data92 (.PAD(PI_Inst_Cahe_readData_data[92]), .C(WIRE_Inst_Cahe_readData_data[92]));
PDIDGZ PAD_Inst_Cahe_readData_data93 (.PAD(PI_Inst_Cahe_readData_data[93]), .C(WIRE_Inst_Cahe_readData_data[93]));
PDIDGZ PAD_Inst_Cahe_readData_data94 (.PAD(PI_Inst_Cahe_readData_data[94]), .C(WIRE_Inst_Cahe_readData_data[94]));
PDIDGZ PAD_Inst_Cahe_readData_data95 (.PAD(PI_Inst_Cahe_readData_data[95]), .C(WIRE_Inst_Cahe_readData_data[95]));
PDIDGZ PAD_Inst_Cahe_readData_data96 (.PAD(PI_Inst_Cahe_readData_data[96]), .C(WIRE_Inst_Cahe_readData_data[96]));
PDIDGZ PAD_Inst_Cahe_readData_data97 (.PAD(PI_Inst_Cahe_readData_data[97]), .C(WIRE_Inst_Cahe_readData_data[97]));
PDIDGZ PAD_Inst_Cahe_readData_data98 (.PAD(PI_Inst_Cahe_readData_data[98]), .C(WIRE_Inst_Cahe_readData_data[98]));
PDIDGZ PAD_Inst_Cahe_readData_data99 (.PAD(PI_Inst_Cahe_readData_data[99]), .C(WIRE_Inst_Cahe_readData_data[99]));
PDIDGZ PAD_Inst_Cahe_readData_data100 (.PAD(PI_Inst_Cahe_readData_data[100]), .C(WIRE_Inst_Cahe_readData_data[100]));
PDIDGZ PAD_Inst_Cahe_readData_data101 (.PAD(PI_Inst_Cahe_readData_data[101]), .C(WIRE_Inst_Cahe_readData_data[101]));
PDIDGZ PAD_Inst_Cahe_readData_data102 (.PAD(PI_Inst_Cahe_readData_data[102]), .C(WIRE_Inst_Cahe_readData_data[102]));
PDIDGZ PAD_Inst_Cahe_readData_data103 (.PAD(PI_Inst_Cahe_readData_data[103]), .C(WIRE_Inst_Cahe_readData_data[103]));
PDIDGZ PAD_Inst_Cahe_readData_data104 (.PAD(PI_Inst_Cahe_readData_data[104]), .C(WIRE_Inst_Cahe_readData_data[104]));
PDIDGZ PAD_Inst_Cahe_readData_data105 (.PAD(PI_Inst_Cahe_readData_data[105]), .C(WIRE_Inst_Cahe_readData_data[105]));
PDIDGZ PAD_Inst_Cahe_readData_data106 (.PAD(PI_Inst_Cahe_readData_data[106]), .C(WIRE_Inst_Cahe_readData_data[106]));
PDIDGZ PAD_Inst_Cahe_readData_data107 (.PAD(PI_Inst_Cahe_readData_data[107]), .C(WIRE_Inst_Cahe_readData_data[107]));
PDIDGZ PAD_Inst_Cahe_readData_data108 (.PAD(PI_Inst_Cahe_readData_data[108]), .C(WIRE_Inst_Cahe_readData_data[108]));
PDIDGZ PAD_Inst_Cahe_readData_data109 (.PAD(PI_Inst_Cahe_readData_data[109]), .C(WIRE_Inst_Cahe_readData_data[109]));
PDIDGZ PAD_Inst_Cahe_readData_data110 (.PAD(PI_Inst_Cahe_readData_data[110]), .C(WIRE_Inst_Cahe_readData_data[110]));
PDIDGZ PAD_Inst_Cahe_readData_data111 (.PAD(PI_Inst_Cahe_readData_data[111]), .C(WIRE_Inst_Cahe_readData_data[111]));
PDIDGZ PAD_Inst_Cahe_readData_data112 (.PAD(PI_Inst_Cahe_readData_data[112]), .C(WIRE_Inst_Cahe_readData_data[112]));
PDIDGZ PAD_Inst_Cahe_readData_data113 (.PAD(PI_Inst_Cahe_readData_data[113]), .C(WIRE_Inst_Cahe_readData_data[113]));
PDIDGZ PAD_Inst_Cahe_readData_data114 (.PAD(PI_Inst_Cahe_readData_data[114]), .C(WIRE_Inst_Cahe_readData_data[114]));
PDIDGZ PAD_Inst_Cahe_readData_data115 (.PAD(PI_Inst_Cahe_readData_data[115]), .C(WIRE_Inst_Cahe_readData_data[115]));
PDIDGZ PAD_Inst_Cahe_readData_data116 (.PAD(PI_Inst_Cahe_readData_data[116]), .C(WIRE_Inst_Cahe_readData_data[116]));
PDIDGZ PAD_Inst_Cahe_readData_data117 (.PAD(PI_Inst_Cahe_readData_data[117]), .C(WIRE_Inst_Cahe_readData_data[117]));
PDIDGZ PAD_Inst_Cahe_readData_data118 (.PAD(PI_Inst_Cahe_readData_data[118]), .C(WIRE_Inst_Cahe_readData_data[118]));
PDIDGZ PAD_Inst_Cahe_readData_data119 (.PAD(PI_Inst_Cahe_readData_data[119]), .C(WIRE_Inst_Cahe_readData_data[119]));
PDIDGZ PAD_Inst_Cahe_readData_data120 (.PAD(PI_Inst_Cahe_readData_data[120]), .C(WIRE_Inst_Cahe_readData_data[120]));
PDIDGZ PAD_Inst_Cahe_readData_data121 (.PAD(PI_Inst_Cahe_readData_data[121]), .C(WIRE_Inst_Cahe_readData_data[121]));
PDIDGZ PAD_Inst_Cahe_readData_data122 (.PAD(PI_Inst_Cahe_readData_data[122]), .C(WIRE_Inst_Cahe_readData_data[122]));
PDIDGZ PAD_Inst_Cahe_readData_data123 (.PAD(PI_Inst_Cahe_readData_data[123]), .C(WIRE_Inst_Cahe_readData_data[123]));
PDIDGZ PAD_Inst_Cahe_readData_data124 (.PAD(PI_Inst_Cahe_readData_data[124]), .C(WIRE_Inst_Cahe_readData_data[124]));
PDIDGZ PAD_Inst_Cahe_readData_data125 (.PAD(PI_Inst_Cahe_readData_data[125]), .C(WIRE_Inst_Cahe_readData_data[125]));
PDIDGZ PAD_Inst_Cahe_readData_data126 (.PAD(PI_Inst_Cahe_readData_data[126]), .C(WIRE_Inst_Cahe_readData_data[126]));
PDIDGZ PAD_Inst_Cahe_readData_data127 (.PAD(PI_Inst_Cahe_readData_data[127]), .C(WIRE_Inst_Cahe_readData_data[127]));

PDIDGZ PAD_Inst_Cahe_readData_valid   (.PAD(PI_Inst_Cahe_readData_valid), .C(WIRE_Inst_Cahe_readData_valid));
PDIDGZ PAD_Inst_Cahe_writeAddr_ready  (.PAD(PI_Inst_Cahe_writeAddr_ready), .C(WIRE_Inst_Cahe_writeAddr_ready));
PDIDGZ PAD_Inst_Cahe_writeData_ready  (.PAD(PI_Inst_Cahe_writeData_ready), .C(WIRE_Inst_Cahe_writeData_ready));

PDIDGZ PAD_Inst_Cahe_writeResp_msg0 (.PAD(PI_Inst_Cahe_writeResp_msg[0]), .C(WIRE_Inst_Cahe_writeResp_msg[0]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg1 (.PAD(PI_Inst_Cahe_writeResp_msg[1]), .C(WIRE_Inst_Cahe_writeResp_msg[1]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg2 (.PAD(PI_Inst_Cahe_writeResp_msg[2]), .C(WIRE_Inst_Cahe_writeResp_msg[2]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg3 (.PAD(PI_Inst_Cahe_writeResp_msg[3]), .C(WIRE_Inst_Cahe_writeResp_msg[3]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg4 (.PAD(PI_Inst_Cahe_writeResp_msg[4]), .C(WIRE_Inst_Cahe_writeResp_msg[4]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg5 (.PAD(PI_Inst_Cahe_writeResp_msg[5]), .C(WIRE_Inst_Cahe_writeResp_msg[5]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg6 (.PAD(PI_Inst_Cahe_writeResp_msg[6]), .C(WIRE_Inst_Cahe_writeResp_msg[6]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg7 (.PAD(PI_Inst_Cahe_writeResp_msg[7]), .C(WIRE_Inst_Cahe_writeResp_msg[7]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg8 (.PAD(PI_Inst_Cahe_writeResp_msg[8]), .C(WIRE_Inst_Cahe_writeResp_msg[8]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg9 (.PAD(PI_Inst_Cahe_writeResp_msg[9]), .C(WIRE_Inst_Cahe_writeResp_msg[9]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg10 (.PAD(PI_Inst_Cahe_writeResp_msg[10]), .C(WIRE_Inst_Cahe_writeResp_msg[10]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg11 (.PAD(PI_Inst_Cahe_writeResp_msg[11]), .C(WIRE_Inst_Cahe_writeResp_msg[11]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg12 (.PAD(PI_Inst_Cahe_writeResp_msg[12]), .C(WIRE_Inst_Cahe_writeResp_msg[12]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg13 (.PAD(PI_Inst_Cahe_writeResp_msg[13]), .C(WIRE_Inst_Cahe_writeResp_msg[13]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg14 (.PAD(PI_Inst_Cahe_writeResp_msg[14]), .C(WIRE_Inst_Cahe_writeResp_msg[14]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg15 (.PAD(PI_Inst_Cahe_writeResp_msg[15]), .C(WIRE_Inst_Cahe_writeResp_msg[15]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg16 (.PAD(PI_Inst_Cahe_writeResp_msg[16]), .C(WIRE_Inst_Cahe_writeResp_msg[16]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg17 (.PAD(PI_Inst_Cahe_writeResp_msg[17]), .C(WIRE_Inst_Cahe_writeResp_msg[17]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg18 (.PAD(PI_Inst_Cahe_writeResp_msg[18]), .C(WIRE_Inst_Cahe_writeResp_msg[18]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg19 (.PAD(PI_Inst_Cahe_writeResp_msg[19]), .C(WIRE_Inst_Cahe_writeResp_msg[19]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg20 (.PAD(PI_Inst_Cahe_writeResp_msg[20]), .C(WIRE_Inst_Cahe_writeResp_msg[20]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg21 (.PAD(PI_Inst_Cahe_writeResp_msg[21]), .C(WIRE_Inst_Cahe_writeResp_msg[21]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg22 (.PAD(PI_Inst_Cahe_writeResp_msg[22]), .C(WIRE_Inst_Cahe_writeResp_msg[22]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg23 (.PAD(PI_Inst_Cahe_writeResp_msg[23]), .C(WIRE_Inst_Cahe_writeResp_msg[23]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg24 (.PAD(PI_Inst_Cahe_writeResp_msg[24]), .C(WIRE_Inst_Cahe_writeResp_msg[24]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg25 (.PAD(PI_Inst_Cahe_writeResp_msg[25]), .C(WIRE_Inst_Cahe_writeResp_msg[25]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg26 (.PAD(PI_Inst_Cahe_writeResp_msg[26]), .C(WIRE_Inst_Cahe_writeResp_msg[26]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg27 (.PAD(PI_Inst_Cahe_writeResp_msg[27]), .C(WIRE_Inst_Cahe_writeResp_msg[27]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg28 (.PAD(PI_Inst_Cahe_writeResp_msg[28]), .C(WIRE_Inst_Cahe_writeResp_msg[28]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg29 (.PAD(PI_Inst_Cahe_writeResp_msg[29]), .C(WIRE_Inst_Cahe_writeResp_msg[29]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg30 (.PAD(PI_Inst_Cahe_writeResp_msg[30]), .C(WIRE_Inst_Cahe_writeResp_msg[30]));
PDIDGZ PAD_Inst_Cahe_writeResp_msg31 (.PAD(PI_Inst_Cahe_writeResp_msg[31]), .C(WIRE_Inst_Cahe_writeResp_msg[31]));

PDIDGZ PAD_Inst_Cahe_writeResp_valid  (.PAD(PI_Inst_Cahe_writeResp_valid), .C(WIRE_Inst_Cahe_writeResp_valid));
PDIDGZ PAD_clk (.PAD(PI_clk), .C(WIRE_clk));
PDIDGZ PAD_rst (.PAD(PI_rst), .C(WIRE_rst));

// CORNER2
PDIDGZ PAD_Data_Cahe_readAddr_ready  (.PAD(PI_Data_Cahe_readAddr_ready), .C(WIRE_Data_Cahe_readAddr_ready));

PDIDGZ PAD_Data_Cahe_readData_data0 (.PAD(PI_Data_Cahe_readData_data[0]), .C(WIRE_Data_Cahe_readData_data[0]));
PDIDGZ PAD_Data_Cahe_readData_data1 (.PAD(PI_Data_Cahe_readData_data[1]), .C(WIRE_Data_Cahe_readData_data[1]));
PDIDGZ PAD_Data_Cahe_readData_data2 (.PAD(PI_Data_Cahe_readData_data[2]), .C(WIRE_Data_Cahe_readData_data[2]));
PDIDGZ PAD_Data_Cahe_readData_data3 (.PAD(PI_Data_Cahe_readData_data[3]), .C(WIRE_Data_Cahe_readData_data[3]));
PDIDGZ PAD_Data_Cahe_readData_data4 (.PAD(PI_Data_Cahe_readData_data[4]), .C(WIRE_Data_Cahe_readData_data[4]));
PDIDGZ PAD_Data_Cahe_readData_data5 (.PAD(PI_Data_Cahe_readData_data[5]), .C(WIRE_Data_Cahe_readData_data[5]));
PDIDGZ PAD_Data_Cahe_readData_data6 (.PAD(PI_Data_Cahe_readData_data[6]), .C(WIRE_Data_Cahe_readData_data[6]));
PDIDGZ PAD_Data_Cahe_readData_data7 (.PAD(PI_Data_Cahe_readData_data[7]), .C(WIRE_Data_Cahe_readData_data[7]));
PDIDGZ PAD_Data_Cahe_readData_data8 (.PAD(PI_Data_Cahe_readData_data[8]), .C(WIRE_Data_Cahe_readData_data[8]));
PDIDGZ PAD_Data_Cahe_readData_data9 (.PAD(PI_Data_Cahe_readData_data[9]), .C(WIRE_Data_Cahe_readData_data[9]));
PDIDGZ PAD_Data_Cahe_readData_data10 (.PAD(PI_Data_Cahe_readData_data[10]), .C(WIRE_Data_Cahe_readData_data[10]));
PDIDGZ PAD_Data_Cahe_readData_data11 (.PAD(PI_Data_Cahe_readData_data[11]), .C(WIRE_Data_Cahe_readData_data[11]));
PDIDGZ PAD_Data_Cahe_readData_data12 (.PAD(PI_Data_Cahe_readData_data[12]), .C(WIRE_Data_Cahe_readData_data[12]));
PDIDGZ PAD_Data_Cahe_readData_data13 (.PAD(PI_Data_Cahe_readData_data[13]), .C(WIRE_Data_Cahe_readData_data[13]));
PDIDGZ PAD_Data_Cahe_readData_data14 (.PAD(PI_Data_Cahe_readData_data[14]), .C(WIRE_Data_Cahe_readData_data[14]));
PDIDGZ PAD_Data_Cahe_readData_data15 (.PAD(PI_Data_Cahe_readData_data[15]), .C(WIRE_Data_Cahe_readData_data[15]));
PDIDGZ PAD_Data_Cahe_readData_data16 (.PAD(PI_Data_Cahe_readData_data[16]), .C(WIRE_Data_Cahe_readData_data[16]));
PDIDGZ PAD_Data_Cahe_readData_data17 (.PAD(PI_Data_Cahe_readData_data[17]), .C(WIRE_Data_Cahe_readData_data[17]));
PDIDGZ PAD_Data_Cahe_readData_data18 (.PAD(PI_Data_Cahe_readData_data[18]), .C(WIRE_Data_Cahe_readData_data[18]));
PDIDGZ PAD_Data_Cahe_readData_data19 (.PAD(PI_Data_Cahe_readData_data[19]), .C(WIRE_Data_Cahe_readData_data[19]));
PDIDGZ PAD_Data_Cahe_readData_data20 (.PAD(PI_Data_Cahe_readData_data[20]), .C(WIRE_Data_Cahe_readData_data[20]));
PDIDGZ PAD_Data_Cahe_readData_data21 (.PAD(PI_Data_Cahe_readData_data[21]), .C(WIRE_Data_Cahe_readData_data[21]));
PDIDGZ PAD_Data_Cahe_readData_data22 (.PAD(PI_Data_Cahe_readData_data[22]), .C(WIRE_Data_Cahe_readData_data[22]));
PDIDGZ PAD_Data_Cahe_readData_data23 (.PAD(PI_Data_Cahe_readData_data[23]), .C(WIRE_Data_Cahe_readData_data[23]));
PDIDGZ PAD_Data_Cahe_readData_data24 (.PAD(PI_Data_Cahe_readData_data[24]), .C(WIRE_Data_Cahe_readData_data[24]));
PDIDGZ PAD_Data_Cahe_readData_data25 (.PAD(PI_Data_Cahe_readData_data[25]), .C(WIRE_Data_Cahe_readData_data[25]));
PDIDGZ PAD_Data_Cahe_readData_data26 (.PAD(PI_Data_Cahe_readData_data[26]), .C(WIRE_Data_Cahe_readData_data[26]));
PDIDGZ PAD_Data_Cahe_readData_data27 (.PAD(PI_Data_Cahe_readData_data[27]), .C(WIRE_Data_Cahe_readData_data[27]));
PDIDGZ PAD_Data_Cahe_readData_data28 (.PAD(PI_Data_Cahe_readData_data[28]), .C(WIRE_Data_Cahe_readData_data[28]));
PDIDGZ PAD_Data_Cahe_readData_data29 (.PAD(PI_Data_Cahe_readData_data[29]), .C(WIRE_Data_Cahe_readData_data[29]));
PDIDGZ PAD_Data_Cahe_readData_data30 (.PAD(PI_Data_Cahe_readData_data[30]), .C(WIRE_Data_Cahe_readData_data[30]));
PDIDGZ PAD_Data_Cahe_readData_data31 (.PAD(PI_Data_Cahe_readData_data[31]), .C(WIRE_Data_Cahe_readData_data[31]));
PDIDGZ PAD_Data_Cahe_readData_data32 (.PAD(PI_Data_Cahe_readData_data[32]), .C(WIRE_Data_Cahe_readData_data[32]));
PDIDGZ PAD_Data_Cahe_readData_data33 (.PAD(PI_Data_Cahe_readData_data[33]), .C(WIRE_Data_Cahe_readData_data[33]));
PDIDGZ PAD_Data_Cahe_readData_data34 (.PAD(PI_Data_Cahe_readData_data[34]), .C(WIRE_Data_Cahe_readData_data[34]));
PDIDGZ PAD_Data_Cahe_readData_data35 (.PAD(PI_Data_Cahe_readData_data[35]), .C(WIRE_Data_Cahe_readData_data[35]));
PDIDGZ PAD_Data_Cahe_readData_data36 (.PAD(PI_Data_Cahe_readData_data[36]), .C(WIRE_Data_Cahe_readData_data[36]));
PDIDGZ PAD_Data_Cahe_readData_data37 (.PAD(PI_Data_Cahe_readData_data[37]), .C(WIRE_Data_Cahe_readData_data[37]));
PDIDGZ PAD_Data_Cahe_readData_data38 (.PAD(PI_Data_Cahe_readData_data[38]), .C(WIRE_Data_Cahe_readData_data[38]));
PDIDGZ PAD_Data_Cahe_readData_data39 (.PAD(PI_Data_Cahe_readData_data[39]), .C(WIRE_Data_Cahe_readData_data[39]));
PDIDGZ PAD_Data_Cahe_readData_data40 (.PAD(PI_Data_Cahe_readData_data[40]), .C(WIRE_Data_Cahe_readData_data[40]));
PDIDGZ PAD_Data_Cahe_readData_data41 (.PAD(PI_Data_Cahe_readData_data[41]), .C(WIRE_Data_Cahe_readData_data[41]));
PDIDGZ PAD_Data_Cahe_readData_data42 (.PAD(PI_Data_Cahe_readData_data[42]), .C(WIRE_Data_Cahe_readData_data[42]));
PDIDGZ PAD_Data_Cahe_readData_data43 (.PAD(PI_Data_Cahe_readData_data[43]), .C(WIRE_Data_Cahe_readData_data[43]));
PDIDGZ PAD_Data_Cahe_readData_data44 (.PAD(PI_Data_Cahe_readData_data[44]), .C(WIRE_Data_Cahe_readData_data[44]));
PDIDGZ PAD_Data_Cahe_readData_data45 (.PAD(PI_Data_Cahe_readData_data[45]), .C(WIRE_Data_Cahe_readData_data[45]));
PDIDGZ PAD_Data_Cahe_readData_data46 (.PAD(PI_Data_Cahe_readData_data[46]), .C(WIRE_Data_Cahe_readData_data[46]));
PDIDGZ PAD_Data_Cahe_readData_data47 (.PAD(PI_Data_Cahe_readData_data[47]), .C(WIRE_Data_Cahe_readData_data[47]));
PDIDGZ PAD_Data_Cahe_readData_data48 (.PAD(PI_Data_Cahe_readData_data[48]), .C(WIRE_Data_Cahe_readData_data[48]));
PDIDGZ PAD_Data_Cahe_readData_data49 (.PAD(PI_Data_Cahe_readData_data[49]), .C(WIRE_Data_Cahe_readData_data[49]));
PDIDGZ PAD_Data_Cahe_readData_data50 (.PAD(PI_Data_Cahe_readData_data[50]), .C(WIRE_Data_Cahe_readData_data[50]));
PDIDGZ PAD_Data_Cahe_readData_data51 (.PAD(PI_Data_Cahe_readData_data[51]), .C(WIRE_Data_Cahe_readData_data[51]));
PDIDGZ PAD_Data_Cahe_readData_data52 (.PAD(PI_Data_Cahe_readData_data[52]), .C(WIRE_Data_Cahe_readData_data[52]));
PDIDGZ PAD_Data_Cahe_readData_data53 (.PAD(PI_Data_Cahe_readData_data[53]), .C(WIRE_Data_Cahe_readData_data[53]));
PDIDGZ PAD_Data_Cahe_readData_data54 (.PAD(PI_Data_Cahe_readData_data[54]), .C(WIRE_Data_Cahe_readData_data[54]));
PDIDGZ PAD_Data_Cahe_readData_data55 (.PAD(PI_Data_Cahe_readData_data[55]), .C(WIRE_Data_Cahe_readData_data[55]));
PDIDGZ PAD_Data_Cahe_readData_data56 (.PAD(PI_Data_Cahe_readData_data[56]), .C(WIRE_Data_Cahe_readData_data[56]));
PDIDGZ PAD_Data_Cahe_readData_data57 (.PAD(PI_Data_Cahe_readData_data[57]), .C(WIRE_Data_Cahe_readData_data[57]));
PDIDGZ PAD_Data_Cahe_readData_data58 (.PAD(PI_Data_Cahe_readData_data[58]), .C(WIRE_Data_Cahe_readData_data[58]));
PDIDGZ PAD_Data_Cahe_readData_data59 (.PAD(PI_Data_Cahe_readData_data[59]), .C(WIRE_Data_Cahe_readData_data[59]));
PDIDGZ PAD_Data_Cahe_readData_data60 (.PAD(PI_Data_Cahe_readData_data[60]), .C(WIRE_Data_Cahe_readData_data[60]));
PDIDGZ PAD_Data_Cahe_readData_data61 (.PAD(PI_Data_Cahe_readData_data[61]), .C(WIRE_Data_Cahe_readData_data[61]));
PDIDGZ PAD_Data_Cahe_readData_data62 (.PAD(PI_Data_Cahe_readData_data[62]), .C(WIRE_Data_Cahe_readData_data[62]));
PDIDGZ PAD_Data_Cahe_readData_data63 (.PAD(PI_Data_Cahe_readData_data[63]), .C(WIRE_Data_Cahe_readData_data[63]));
PDIDGZ PAD_Data_Cahe_readData_data64 (.PAD(PI_Data_Cahe_readData_data[64]), .C(WIRE_Data_Cahe_readData_data[64]));
PDIDGZ PAD_Data_Cahe_readData_data65 (.PAD(PI_Data_Cahe_readData_data[65]), .C(WIRE_Data_Cahe_readData_data[65]));
PDIDGZ PAD_Data_Cahe_readData_data66 (.PAD(PI_Data_Cahe_readData_data[66]), .C(WIRE_Data_Cahe_readData_data[66]));
PDIDGZ PAD_Data_Cahe_readData_data67 (.PAD(PI_Data_Cahe_readData_data[67]), .C(WIRE_Data_Cahe_readData_data[67]));
PDIDGZ PAD_Data_Cahe_readData_data68 (.PAD(PI_Data_Cahe_readData_data[68]), .C(WIRE_Data_Cahe_readData_data[68]));
PDIDGZ PAD_Data_Cahe_readData_data69 (.PAD(PI_Data_Cahe_readData_data[69]), .C(WIRE_Data_Cahe_readData_data[69]));
PDIDGZ PAD_Data_Cahe_readData_data70 (.PAD(PI_Data_Cahe_readData_data[70]), .C(WIRE_Data_Cahe_readData_data[70]));
PDIDGZ PAD_Data_Cahe_readData_data71 (.PAD(PI_Data_Cahe_readData_data[71]), .C(WIRE_Data_Cahe_readData_data[71]));
PDIDGZ PAD_Data_Cahe_readData_data72 (.PAD(PI_Data_Cahe_readData_data[72]), .C(WIRE_Data_Cahe_readData_data[72]));
PDIDGZ PAD_Data_Cahe_readData_data73 (.PAD(PI_Data_Cahe_readData_data[73]), .C(WIRE_Data_Cahe_readData_data[73]));
PDIDGZ PAD_Data_Cahe_readData_data74 (.PAD(PI_Data_Cahe_readData_data[74]), .C(WIRE_Data_Cahe_readData_data[74]));
PDIDGZ PAD_Data_Cahe_readData_data75 (.PAD(PI_Data_Cahe_readData_data[75]), .C(WIRE_Data_Cahe_readData_data[75]));
PDIDGZ PAD_Data_Cahe_readData_data76 (.PAD(PI_Data_Cahe_readData_data[76]), .C(WIRE_Data_Cahe_readData_data[76]));
PDIDGZ PAD_Data_Cahe_readData_data77 (.PAD(PI_Data_Cahe_readData_data[77]), .C(WIRE_Data_Cahe_readData_data[77]));
PDIDGZ PAD_Data_Cahe_readData_data78 (.PAD(PI_Data_Cahe_readData_data[78]), .C(WIRE_Data_Cahe_readData_data[78]));
PDIDGZ PAD_Data_Cahe_readData_data79 (.PAD(PI_Data_Cahe_readData_data[79]), .C(WIRE_Data_Cahe_readData_data[79]));
PDIDGZ PAD_Data_Cahe_readData_data80 (.PAD(PI_Data_Cahe_readData_data[80]), .C(WIRE_Data_Cahe_readData_data[80]));
PDIDGZ PAD_Data_Cahe_readData_data81 (.PAD(PI_Data_Cahe_readData_data[81]), .C(WIRE_Data_Cahe_readData_data[81]));
PDIDGZ PAD_Data_Cahe_readData_data82 (.PAD(PI_Data_Cahe_readData_data[82]), .C(WIRE_Data_Cahe_readData_data[82]));
PDIDGZ PAD_Data_Cahe_readData_data83 (.PAD(PI_Data_Cahe_readData_data[83]), .C(WIRE_Data_Cahe_readData_data[83]));
PDIDGZ PAD_Data_Cahe_readData_data84 (.PAD(PI_Data_Cahe_readData_data[84]), .C(WIRE_Data_Cahe_readData_data[84]));
PDIDGZ PAD_Data_Cahe_readData_data85 (.PAD(PI_Data_Cahe_readData_data[85]), .C(WIRE_Data_Cahe_readData_data[85]));
PDIDGZ PAD_Data_Cahe_readData_data86 (.PAD(PI_Data_Cahe_readData_data[86]), .C(WIRE_Data_Cahe_readData_data[86]));
PDIDGZ PAD_Data_Cahe_readData_data87 (.PAD(PI_Data_Cahe_readData_data[87]), .C(WIRE_Data_Cahe_readData_data[87]));
PDIDGZ PAD_Data_Cahe_readData_data88 (.PAD(PI_Data_Cahe_readData_data[88]), .C(WIRE_Data_Cahe_readData_data[88]));
PDIDGZ PAD_Data_Cahe_readData_data89 (.PAD(PI_Data_Cahe_readData_data[89]), .C(WIRE_Data_Cahe_readData_data[89]));
PDIDGZ PAD_Data_Cahe_readData_data90 (.PAD(PI_Data_Cahe_readData_data[90]), .C(WIRE_Data_Cahe_readData_data[90]));
PDIDGZ PAD_Data_Cahe_readData_data91 (.PAD(PI_Data_Cahe_readData_data[91]), .C(WIRE_Data_Cahe_readData_data[91]));
PDIDGZ PAD_Data_Cahe_readData_data92 (.PAD(PI_Data_Cahe_readData_data[92]), .C(WIRE_Data_Cahe_readData_data[92]));
PDIDGZ PAD_Data_Cahe_readData_data93 (.PAD(PI_Data_Cahe_readData_data[93]), .C(WIRE_Data_Cahe_readData_data[93]));
PDIDGZ PAD_Data_Cahe_readData_data94 (.PAD(PI_Data_Cahe_readData_data[94]), .C(WIRE_Data_Cahe_readData_data[94]));
PDIDGZ PAD_Data_Cahe_readData_data95 (.PAD(PI_Data_Cahe_readData_data[95]), .C(WIRE_Data_Cahe_readData_data[95]));
PDIDGZ PAD_Data_Cahe_readData_data96 (.PAD(PI_Data_Cahe_readData_data[96]), .C(WIRE_Data_Cahe_readData_data[96]));
PDIDGZ PAD_Data_Cahe_readData_data97 (.PAD(PI_Data_Cahe_readData_data[97]), .C(WIRE_Data_Cahe_readData_data[97]));
PDIDGZ PAD_Data_Cahe_readData_data98 (.PAD(PI_Data_Cahe_readData_data[98]), .C(WIRE_Data_Cahe_readData_data[98]));
PDIDGZ PAD_Data_Cahe_readData_data99 (.PAD(PI_Data_Cahe_readData_data[99]), .C(WIRE_Data_Cahe_readData_data[99]));
PDIDGZ PAD_Data_Cahe_readData_data100 (.PAD(PI_Data_Cahe_readData_data[100]), .C(WIRE_Data_Cahe_readData_data[100]));
PDIDGZ PAD_Data_Cahe_readData_data101 (.PAD(PI_Data_Cahe_readData_data[101]), .C(WIRE_Data_Cahe_readData_data[101]));
PDIDGZ PAD_Data_Cahe_readData_data102 (.PAD(PI_Data_Cahe_readData_data[102]), .C(WIRE_Data_Cahe_readData_data[102]));
PDIDGZ PAD_Data_Cahe_readData_data103 (.PAD(PI_Data_Cahe_readData_data[103]), .C(WIRE_Data_Cahe_readData_data[103]));
PDIDGZ PAD_Data_Cahe_readData_data104 (.PAD(PI_Data_Cahe_readData_data[104]), .C(WIRE_Data_Cahe_readData_data[104]));
PDIDGZ PAD_Data_Cahe_readData_data105 (.PAD(PI_Data_Cahe_readData_data[105]), .C(WIRE_Data_Cahe_readData_data[105]));
PDIDGZ PAD_Data_Cahe_readData_data106 (.PAD(PI_Data_Cahe_readData_data[106]), .C(WIRE_Data_Cahe_readData_data[106]));
PDIDGZ PAD_Data_Cahe_readData_data107 (.PAD(PI_Data_Cahe_readData_data[107]), .C(WIRE_Data_Cahe_readData_data[107]));
PDIDGZ PAD_Data_Cahe_readData_data108 (.PAD(PI_Data_Cahe_readData_data[108]), .C(WIRE_Data_Cahe_readData_data[108]));
PDIDGZ PAD_Data_Cahe_readData_data109 (.PAD(PI_Data_Cahe_readData_data[109]), .C(WIRE_Data_Cahe_readData_data[109]));
PDIDGZ PAD_Data_Cahe_readData_data110 (.PAD(PI_Data_Cahe_readData_data[110]), .C(WIRE_Data_Cahe_readData_data[110]));
PDIDGZ PAD_Data_Cahe_readData_data111 (.PAD(PI_Data_Cahe_readData_data[111]), .C(WIRE_Data_Cahe_readData_data[111]));
PDIDGZ PAD_Data_Cahe_readData_data112 (.PAD(PI_Data_Cahe_readData_data[112]), .C(WIRE_Data_Cahe_readData_data[112]));
PDIDGZ PAD_Data_Cahe_readData_data113 (.PAD(PI_Data_Cahe_readData_data[113]), .C(WIRE_Data_Cahe_readData_data[113]));
PDIDGZ PAD_Data_Cahe_readData_data114 (.PAD(PI_Data_Cahe_readData_data[114]), .C(WIRE_Data_Cahe_readData_data[114]));
PDIDGZ PAD_Data_Cahe_readData_data115 (.PAD(PI_Data_Cahe_readData_data[115]), .C(WIRE_Data_Cahe_readData_data[115]));
PDIDGZ PAD_Data_Cahe_readData_data116 (.PAD(PI_Data_Cahe_readData_data[116]), .C(WIRE_Data_Cahe_readData_data[116]));
PDIDGZ PAD_Data_Cahe_readData_data117 (.PAD(PI_Data_Cahe_readData_data[117]), .C(WIRE_Data_Cahe_readData_data[117]));
PDIDGZ PAD_Data_Cahe_readData_data118 (.PAD(PI_Data_Cahe_readData_data[118]), .C(WIRE_Data_Cahe_readData_data[118]));
PDIDGZ PAD_Data_Cahe_readData_data119 (.PAD(PI_Data_Cahe_readData_data[119]), .C(WIRE_Data_Cahe_readData_data[119]));
PDIDGZ PAD_Data_Cahe_readData_data120 (.PAD(PI_Data_Cahe_readData_data[120]), .C(WIRE_Data_Cahe_readData_data[120]));
PDIDGZ PAD_Data_Cahe_readData_data121 (.PAD(PI_Data_Cahe_readData_data[121]), .C(WIRE_Data_Cahe_readData_data[121]));
PDIDGZ PAD_Data_Cahe_readData_data122 (.PAD(PI_Data_Cahe_readData_data[122]), .C(WIRE_Data_Cahe_readData_data[122]));
PDIDGZ PAD_Data_Cahe_readData_data123 (.PAD(PI_Data_Cahe_readData_data[123]), .C(WIRE_Data_Cahe_readData_data[123]));
PDIDGZ PAD_Data_Cahe_readData_data124 (.PAD(PI_Data_Cahe_readData_data[124]), .C(WIRE_Data_Cahe_readData_data[124]));
PDIDGZ PAD_Data_Cahe_readData_data125 (.PAD(PI_Data_Cahe_readData_data[125]), .C(WIRE_Data_Cahe_readData_data[125]));
PDIDGZ PAD_Data_Cahe_readData_data126 (.PAD(PI_Data_Cahe_readData_data[126]), .C(WIRE_Data_Cahe_readData_data[126]));
PDIDGZ PAD_Data_Cahe_readData_data127 (.PAD(PI_Data_Cahe_readData_data[127]), .C(WIRE_Data_Cahe_readData_data[127]));

PDIDGZ PAD_Data_Cahe_readData_valid  (.PAD(PI_Data_Cahe_readData_valid), .C(WIRE_Data_Cahe_readData_valid));
PDIDGZ PAD_Data_Cahe_writeAddr_ready (.PAD(PI_Data_Cahe_writeAddr_ready), .C(WIRE_Data_Cahe_writeAddr_ready));
PDIDGZ PAD_Data_Cahe_writeData_ready (.PAD(PI_Data_Cahe_writeData_ready), .C(WIRE_Data_Cahe_writeData_ready));

PDIDGZ PAD_Data_Cahe_writeResp_msg0 (.PAD(PI_Data_Cahe_writeResp_msg[0]), .C(WIRE_Data_Cahe_writeResp_msg[0]));
PDIDGZ PAD_Data_Cahe_writeResp_msg1 (.PAD(PI_Data_Cahe_writeResp_msg[1]), .C(WIRE_Data_Cahe_writeResp_msg[1]));
PDIDGZ PAD_Data_Cahe_writeResp_msg2 (.PAD(PI_Data_Cahe_writeResp_msg[2]), .C(WIRE_Data_Cahe_writeResp_msg[2]));
PDIDGZ PAD_Data_Cahe_writeResp_msg3 (.PAD(PI_Data_Cahe_writeResp_msg[3]), .C(WIRE_Data_Cahe_writeResp_msg[3]));
PDIDGZ PAD_Data_Cahe_writeResp_msg4 (.PAD(PI_Data_Cahe_writeResp_msg[4]), .C(WIRE_Data_Cahe_writeResp_msg[4]));
PDIDGZ PAD_Data_Cahe_writeResp_msg5 (.PAD(PI_Data_Cahe_writeResp_msg[5]), .C(WIRE_Data_Cahe_writeResp_msg[5]));
PDIDGZ PAD_Data_Cahe_writeResp_msg6 (.PAD(PI_Data_Cahe_writeResp_msg[6]), .C(WIRE_Data_Cahe_writeResp_msg[6]));
PDIDGZ PAD_Data_Cahe_writeResp_msg7 (.PAD(PI_Data_Cahe_writeResp_msg[7]), .C(WIRE_Data_Cahe_writeResp_msg[7]));
PDIDGZ PAD_Data_Cahe_writeResp_msg8 (.PAD(PI_Data_Cahe_writeResp_msg[8]), .C(WIRE_Data_Cahe_writeResp_msg[8]));
PDIDGZ PAD_Data_Cahe_writeResp_msg9 (.PAD(PI_Data_Cahe_writeResp_msg[9]), .C(WIRE_Data_Cahe_writeResp_msg[9]));
PDIDGZ PAD_Data_Cahe_writeResp_msg10 (.PAD(PI_Data_Cahe_writeResp_msg[10]), .C(WIRE_Data_Cahe_writeResp_msg[10]));
PDIDGZ PAD_Data_Cahe_writeResp_msg11 (.PAD(PI_Data_Cahe_writeResp_msg[11]), .C(WIRE_Data_Cahe_writeResp_msg[11]));
PDIDGZ PAD_Data_Cahe_writeResp_msg12 (.PAD(PI_Data_Cahe_writeResp_msg[12]), .C(WIRE_Data_Cahe_writeResp_msg[12]));
PDIDGZ PAD_Data_Cahe_writeResp_msg13 (.PAD(PI_Data_Cahe_writeResp_msg[13]), .C(WIRE_Data_Cahe_writeResp_msg[13]));
PDIDGZ PAD_Data_Cahe_writeResp_msg14 (.PAD(PI_Data_Cahe_writeResp_msg[14]), .C(WIRE_Data_Cahe_writeResp_msg[14]));
PDIDGZ PAD_Data_Cahe_writeResp_msg15 (.PAD(PI_Data_Cahe_writeResp_msg[15]), .C(WIRE_Data_Cahe_writeResp_msg[15]));
PDIDGZ PAD_Data_Cahe_writeResp_msg16 (.PAD(PI_Data_Cahe_writeResp_msg[16]), .C(WIRE_Data_Cahe_writeResp_msg[16]));
PDIDGZ PAD_Data_Cahe_writeResp_msg17 (.PAD(PI_Data_Cahe_writeResp_msg[17]), .C(WIRE_Data_Cahe_writeResp_msg[17]));
PDIDGZ PAD_Data_Cahe_writeResp_msg18 (.PAD(PI_Data_Cahe_writeResp_msg[18]), .C(WIRE_Data_Cahe_writeResp_msg[18]));
PDIDGZ PAD_Data_Cahe_writeResp_msg19 (.PAD(PI_Data_Cahe_writeResp_msg[19]), .C(WIRE_Data_Cahe_writeResp_msg[19]));
PDIDGZ PAD_Data_Cahe_writeResp_msg20 (.PAD(PI_Data_Cahe_writeResp_msg[20]), .C(WIRE_Data_Cahe_writeResp_msg[20]));
PDIDGZ PAD_Data_Cahe_writeResp_msg21 (.PAD(PI_Data_Cahe_writeResp_msg[21]), .C(WIRE_Data_Cahe_writeResp_msg[21]));
PDIDGZ PAD_Data_Cahe_writeResp_msg22 (.PAD(PI_Data_Cahe_writeResp_msg[22]), .C(WIRE_Data_Cahe_writeResp_msg[22]));
PDIDGZ PAD_Data_Cahe_writeResp_msg23 (.PAD(PI_Data_Cahe_writeResp_msg[23]), .C(WIRE_Data_Cahe_writeResp_msg[23]));
PDIDGZ PAD_Data_Cahe_writeResp_msg24 (.PAD(PI_Data_Cahe_writeResp_msg[24]), .C(WIRE_Data_Cahe_writeResp_msg[24]));
PDIDGZ PAD_Data_Cahe_writeResp_msg25 (.PAD(PI_Data_Cahe_writeResp_msg[25]), .C(WIRE_Data_Cahe_writeResp_msg[25]));
PDIDGZ PAD_Data_Cahe_writeResp_msg26 (.PAD(PI_Data_Cahe_writeResp_msg[26]), .C(WIRE_Data_Cahe_writeResp_msg[26]));
PDIDGZ PAD_Data_Cahe_writeResp_msg27 (.PAD(PI_Data_Cahe_writeResp_msg[27]), .C(WIRE_Data_Cahe_writeResp_msg[27]));
PDIDGZ PAD_Data_Cahe_writeResp_msg28 (.PAD(PI_Data_Cahe_writeResp_msg[28]), .C(WIRE_Data_Cahe_writeResp_msg[28]));
PDIDGZ PAD_Data_Cahe_writeResp_msg29 (.PAD(PI_Data_Cahe_writeResp_msg[29]), .C(WIRE_Data_Cahe_writeResp_msg[29]));
PDIDGZ PAD_Data_Cahe_writeResp_msg30 (.PAD(PI_Data_Cahe_writeResp_msg[30]), .C(WIRE_Data_Cahe_writeResp_msg[30]));
PDIDGZ PAD_Data_Cahe_writeResp_msg31 (.PAD(PI_Data_Cahe_writeResp_msg[31]), .C(WIRE_Data_Cahe_writeResp_msg[31]));

PDIDGZ PAD_Data_Cahe_writeResp_valid (.PAD(PI_Data_Cahe_writeResp_valid), .C(WIRE_Data_Cahe_writeResp_valid));

// output pads: PDO02CDG (.I(WIRE), .PAD(PO))
// CORNER0
PDIDGZ PAD_halt (.I(WIRE_halt), .C(PO_halt));

// CORNER1
PDO02CDG PAD_Inst_Cahe_readAddr_addr0 (.I(WIRE_Inst_Cahe_readAddr_addr[0]), .PAD(PO_Inst_Cahe_readAddr_addr[0]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr1 (.I(WIRE_Inst_Cahe_readAddr_addr[1]), .PAD(PO_Inst_Cahe_readAddr_addr[1]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr2 (.I(WIRE_Inst_Cahe_readAddr_addr[2]), .PAD(PO_Inst_Cahe_readAddr_addr[2]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr3 (.I(WIRE_Inst_Cahe_readAddr_addr[3]), .PAD(PO_Inst_Cahe_readAddr_addr[3]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr4 (.I(WIRE_Inst_Cahe_readAddr_addr[4]), .PAD(PO_Inst_Cahe_readAddr_addr[4]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr5 (.I(WIRE_Inst_Cahe_readAddr_addr[5]), .PAD(PO_Inst_Cahe_readAddr_addr[5]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr6 (.I(WIRE_Inst_Cahe_readAddr_addr[6]), .PAD(PO_Inst_Cahe_readAddr_addr[6]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr7 (.I(WIRE_Inst_Cahe_readAddr_addr[7]), .PAD(PO_Inst_Cahe_readAddr_addr[7]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr8 (.I(WIRE_Inst_Cahe_readAddr_addr[8]), .PAD(PO_Inst_Cahe_readAddr_addr[8]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr9 (.I(WIRE_Inst_Cahe_readAddr_addr[9]), .PAD(PO_Inst_Cahe_readAddr_addr[9]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr10 (.I(WIRE_Inst_Cahe_readAddr_addr[10]), .PAD(PO_Inst_Cahe_readAddr_addr[10]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr11 (.I(WIRE_Inst_Cahe_readAddr_addr[11]), .PAD(PO_Inst_Cahe_readAddr_addr[11]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr12 (.I(WIRE_Inst_Cahe_readAddr_addr[12]), .PAD(PO_Inst_Cahe_readAddr_addr[12]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr13 (.I(WIRE_Inst_Cahe_readAddr_addr[13]), .PAD(PO_Inst_Cahe_readAddr_addr[13]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr14 (.I(WIRE_Inst_Cahe_readAddr_addr[14]), .PAD(PO_Inst_Cahe_readAddr_addr[14]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr15 (.I(WIRE_Inst_Cahe_readAddr_addr[15]), .PAD(PO_Inst_Cahe_readAddr_addr[15]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr16 (.I(WIRE_Inst_Cahe_readAddr_addr[16]), .PAD(PO_Inst_Cahe_readAddr_addr[16]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr17 (.I(WIRE_Inst_Cahe_readAddr_addr[17]), .PAD(PO_Inst_Cahe_readAddr_addr[17]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr18 (.I(WIRE_Inst_Cahe_readAddr_addr[18]), .PAD(PO_Inst_Cahe_readAddr_addr[18]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr19 (.I(WIRE_Inst_Cahe_readAddr_addr[19]), .PAD(PO_Inst_Cahe_readAddr_addr[19]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr20 (.I(WIRE_Inst_Cahe_readAddr_addr[20]), .PAD(PO_Inst_Cahe_readAddr_addr[20]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr21 (.I(WIRE_Inst_Cahe_readAddr_addr[21]), .PAD(PO_Inst_Cahe_readAddr_addr[21]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr22 (.I(WIRE_Inst_Cahe_readAddr_addr[22]), .PAD(PO_Inst_Cahe_readAddr_addr[22]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr23 (.I(WIRE_Inst_Cahe_readAddr_addr[23]), .PAD(PO_Inst_Cahe_readAddr_addr[23]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr24 (.I(WIRE_Inst_Cahe_readAddr_addr[24]), .PAD(PO_Inst_Cahe_readAddr_addr[24]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr25 (.I(WIRE_Inst_Cahe_readAddr_addr[25]), .PAD(PO_Inst_Cahe_readAddr_addr[25]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr26 (.I(WIRE_Inst_Cahe_readAddr_addr[26]), .PAD(PO_Inst_Cahe_readAddr_addr[26]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr27 (.I(WIRE_Inst_Cahe_readAddr_addr[27]), .PAD(PO_Inst_Cahe_readAddr_addr[27]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr28 (.I(WIRE_Inst_Cahe_readAddr_addr[28]), .PAD(PO_Inst_Cahe_readAddr_addr[28]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr29 (.I(WIRE_Inst_Cahe_readAddr_addr[29]), .PAD(PO_Inst_Cahe_readAddr_addr[29]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr30 (.I(WIRE_Inst_Cahe_readAddr_addr[30]), .PAD(PO_Inst_Cahe_readAddr_addr[30]));
PDO02CDG PAD_Inst_Cahe_readAddr_addr31 (.I(WIRE_Inst_Cahe_readAddr_addr[31]), .PAD(PO_Inst_Cahe_readAddr_addr[31]));

PDO02CDG PAD_Inst_Cahe_readAddr_valid  (.I(WIRE_Inst_Cahe_readAddr_valid), .PAD(PO_Inst_Cahe_readAddr_valid));
PDO02CDG PAD_Inst_Cahe_readData_ready  (.I(WIRE_Inst_Cahe_readData_ready), .PAD(PO_Inst_Cahe_readData_ready));

PDO02CDG PAD_Inst_Cahe_writeAddr_addr0 (.I(WIRE_Inst_Cahe_writeAddr_addr[0]), .PAD(PO_Inst_Cahe_writeAddr_addr[0]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr1 (.I(WIRE_Inst_Cahe_writeAddr_addr[1]), .PAD(PO_Inst_Cahe_writeAddr_addr[1]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr2 (.I(WIRE_Inst_Cahe_writeAddr_addr[2]), .PAD(PO_Inst_Cahe_writeAddr_addr[2]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr3 (.I(WIRE_Inst_Cahe_writeAddr_addr[3]), .PAD(PO_Inst_Cahe_writeAddr_addr[3]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr4 (.I(WIRE_Inst_Cahe_writeAddr_addr[4]), .PAD(PO_Inst_Cahe_writeAddr_addr[4]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr5 (.I(WIRE_Inst_Cahe_writeAddr_addr[5]), .PAD(PO_Inst_Cahe_writeAddr_addr[5]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr6 (.I(WIRE_Inst_Cahe_writeAddr_addr[6]), .PAD(PO_Inst_Cahe_writeAddr_addr[6]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr7 (.I(WIRE_Inst_Cahe_writeAddr_addr[7]), .PAD(PO_Inst_Cahe_writeAddr_addr[7]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr8 (.I(WIRE_Inst_Cahe_writeAddr_addr[8]), .PAD(PO_Inst_Cahe_writeAddr_addr[8]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr9 (.I(WIRE_Inst_Cahe_writeAddr_addr[9]), .PAD(PO_Inst_Cahe_writeAddr_addr[9]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr10 (.I(WIRE_Inst_Cahe_writeAddr_addr[10]), .PAD(PO_Inst_Cahe_writeAddr_addr[10]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr11 (.I(WIRE_Inst_Cahe_writeAddr_addr[11]), .PAD(PO_Inst_Cahe_writeAddr_addr[11]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr12 (.I(WIRE_Inst_Cahe_writeAddr_addr[12]), .PAD(PO_Inst_Cahe_writeAddr_addr[12]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr13 (.I(WIRE_Inst_Cahe_writeAddr_addr[13]), .PAD(PO_Inst_Cahe_writeAddr_addr[13]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr14 (.I(WIRE_Inst_Cahe_writeAddr_addr[14]), .PAD(PO_Inst_Cahe_writeAddr_addr[14]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr15 (.I(WIRE_Inst_Cahe_writeAddr_addr[15]), .PAD(PO_Inst_Cahe_writeAddr_addr[15]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr16 (.I(WIRE_Inst_Cahe_writeAddr_addr[16]), .PAD(PO_Inst_Cahe_writeAddr_addr[16]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr17 (.I(WIRE_Inst_Cahe_writeAddr_addr[17]), .PAD(PO_Inst_Cahe_writeAddr_addr[17]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr18 (.I(WIRE_Inst_Cahe_writeAddr_addr[18]), .PAD(PO_Inst_Cahe_writeAddr_addr[18]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr19 (.I(WIRE_Inst_Cahe_writeAddr_addr[19]), .PAD(PO_Inst_Cahe_writeAddr_addr[19]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr20 (.I(WIRE_Inst_Cahe_writeAddr_addr[20]), .PAD(PO_Inst_Cahe_writeAddr_addr[20]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr21 (.I(WIRE_Inst_Cahe_writeAddr_addr[21]), .PAD(PO_Inst_Cahe_writeAddr_addr[21]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr22 (.I(WIRE_Inst_Cahe_writeAddr_addr[22]), .PAD(PO_Inst_Cahe_writeAddr_addr[22]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr23 (.I(WIRE_Inst_Cahe_writeAddr_addr[23]), .PAD(PO_Inst_Cahe_writeAddr_addr[23]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr24 (.I(WIRE_Inst_Cahe_writeAddr_addr[24]), .PAD(PO_Inst_Cahe_writeAddr_addr[24]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr25 (.I(WIRE_Inst_Cahe_writeAddr_addr[25]), .PAD(PO_Inst_Cahe_writeAddr_addr[25]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr26 (.I(WIRE_Inst_Cahe_writeAddr_addr[26]), .PAD(PO_Inst_Cahe_writeAddr_addr[26]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr27 (.I(WIRE_Inst_Cahe_writeAddr_addr[27]), .PAD(PO_Inst_Cahe_writeAddr_addr[27]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr28 (.I(WIRE_Inst_Cahe_writeAddr_addr[28]), .PAD(PO_Inst_Cahe_writeAddr_addr[28]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr29 (.I(WIRE_Inst_Cahe_writeAddr_addr[29]), .PAD(PO_Inst_Cahe_writeAddr_addr[29]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr30 (.I(WIRE_Inst_Cahe_writeAddr_addr[30]), .PAD(PO_Inst_Cahe_writeAddr_addr[30]));
PDO02CDG PAD_Inst_Cahe_writeAddr_addr31 (.I(WIRE_Inst_Cahe_writeAddr_addr[31]), .PAD(PO_Inst_Cahe_writeAddr_addr[31]));

PDO02CDG PAD_Inst_Cahe_writeAddr_valid (.I(WIRE_Inst_Cahe_writeAddr_valid), .PAD(PO_Inst_Cahe_writeAddr_valid));

PDO02CDG PAD_Inst_Cahe_writeData_data0 (.I(WIRE_Inst_Cahe_writeData_data[0]), .PAD(PO_Inst_Cahe_writeData_data[0]));
PDO02CDG PAD_Inst_Cahe_writeData_data1 (.I(WIRE_Inst_Cahe_writeData_data[1]), .PAD(PO_Inst_Cahe_writeData_data[1]));
PDO02CDG PAD_Inst_Cahe_writeData_data2 (.I(WIRE_Inst_Cahe_writeData_data[2]), .PAD(PO_Inst_Cahe_writeData_data[2]));
PDO02CDG PAD_Inst_Cahe_writeData_data3 (.I(WIRE_Inst_Cahe_writeData_data[3]), .PAD(PO_Inst_Cahe_writeData_data[3]));
PDO02CDG PAD_Inst_Cahe_writeData_data4 (.I(WIRE_Inst_Cahe_writeData_data[4]), .PAD(PO_Inst_Cahe_writeData_data[4]));
PDO02CDG PAD_Inst_Cahe_writeData_data5 (.I(WIRE_Inst_Cahe_writeData_data[5]), .PAD(PO_Inst_Cahe_writeData_data[5]));
PDO02CDG PAD_Inst_Cahe_writeData_data6 (.I(WIRE_Inst_Cahe_writeData_data[6]), .PAD(PO_Inst_Cahe_writeData_data[6]));
PDO02CDG PAD_Inst_Cahe_writeData_data7 (.I(WIRE_Inst_Cahe_writeData_data[7]), .PAD(PO_Inst_Cahe_writeData_data[7]));
PDO02CDG PAD_Inst_Cahe_writeData_data8 (.I(WIRE_Inst_Cahe_writeData_data[8]), .PAD(PO_Inst_Cahe_writeData_data[8]));
PDO02CDG PAD_Inst_Cahe_writeData_data9 (.I(WIRE_Inst_Cahe_writeData_data[9]), .PAD(PO_Inst_Cahe_writeData_data[9]));
PDO02CDG PAD_Inst_Cahe_writeData_data10 (.I(WIRE_Inst_Cahe_writeData_data[10]), .PAD(PO_Inst_Cahe_writeData_data[10]));
PDO02CDG PAD_Inst_Cahe_writeData_data11 (.I(WIRE_Inst_Cahe_writeData_data[11]), .PAD(PO_Inst_Cahe_writeData_data[11]));
PDO02CDG PAD_Inst_Cahe_writeData_data12 (.I(WIRE_Inst_Cahe_writeData_data[12]), .PAD(PO_Inst_Cahe_writeData_data[12]));
PDO02CDG PAD_Inst_Cahe_writeData_data13 (.I(WIRE_Inst_Cahe_writeData_data[13]), .PAD(PO_Inst_Cahe_writeData_data[13]));
PDO02CDG PAD_Inst_Cahe_writeData_data14 (.I(WIRE_Inst_Cahe_writeData_data[14]), .PAD(PO_Inst_Cahe_writeData_data[14]));
PDO02CDG PAD_Inst_Cahe_writeData_data15 (.I(WIRE_Inst_Cahe_writeData_data[15]), .PAD(PO_Inst_Cahe_writeData_data[15]));
PDO02CDG PAD_Inst_Cahe_writeData_data16 (.I(WIRE_Inst_Cahe_writeData_data[16]), .PAD(PO_Inst_Cahe_writeData_data[16]));
PDO02CDG PAD_Inst_Cahe_writeData_data17 (.I(WIRE_Inst_Cahe_writeData_data[17]), .PAD(PO_Inst_Cahe_writeData_data[17]));
PDO02CDG PAD_Inst_Cahe_writeData_data18 (.I(WIRE_Inst_Cahe_writeData_data[18]), .PAD(PO_Inst_Cahe_writeData_data[18]));
PDO02CDG PAD_Inst_Cahe_writeData_data19 (.I(WIRE_Inst_Cahe_writeData_data[19]), .PAD(PO_Inst_Cahe_writeData_data[19]));
PDO02CDG PAD_Inst_Cahe_writeData_data20 (.I(WIRE_Inst_Cahe_writeData_data[20]), .PAD(PO_Inst_Cahe_writeData_data[20]));
PDO02CDG PAD_Inst_Cahe_writeData_data21 (.I(WIRE_Inst_Cahe_writeData_data[21]), .PAD(PO_Inst_Cahe_writeData_data[21]));
PDO02CDG PAD_Inst_Cahe_writeData_data22 (.I(WIRE_Inst_Cahe_writeData_data[22]), .PAD(PO_Inst_Cahe_writeData_data[22]));
PDO02CDG PAD_Inst_Cahe_writeData_data23 (.I(WIRE_Inst_Cahe_writeData_data[23]), .PAD(PO_Inst_Cahe_writeData_data[23]));
PDO02CDG PAD_Inst_Cahe_writeData_data24 (.I(WIRE_Inst_Cahe_writeData_data[24]), .PAD(PO_Inst_Cahe_writeData_data[24]));
PDO02CDG PAD_Inst_Cahe_writeData_data25 (.I(WIRE_Inst_Cahe_writeData_data[25]), .PAD(PO_Inst_Cahe_writeData_data[25]));
PDO02CDG PAD_Inst_Cahe_writeData_data26 (.I(WIRE_Inst_Cahe_writeData_data[26]), .PAD(PO_Inst_Cahe_writeData_data[26]));
PDO02CDG PAD_Inst_Cahe_writeData_data27 (.I(WIRE_Inst_Cahe_writeData_data[27]), .PAD(PO_Inst_Cahe_writeData_data[27]));
PDO02CDG PAD_Inst_Cahe_writeData_data28 (.I(WIRE_Inst_Cahe_writeData_data[28]), .PAD(PO_Inst_Cahe_writeData_data[28]));
PDO02CDG PAD_Inst_Cahe_writeData_data29 (.I(WIRE_Inst_Cahe_writeData_data[29]), .PAD(PO_Inst_Cahe_writeData_data[29]));
PDO02CDG PAD_Inst_Cahe_writeData_data30 (.I(WIRE_Inst_Cahe_writeData_data[30]), .PAD(PO_Inst_Cahe_writeData_data[30]));
PDO02CDG PAD_Inst_Cahe_writeData_data31 (.I(WIRE_Inst_Cahe_writeData_data[31]), .PAD(PO_Inst_Cahe_writeData_data[31]));
PDO02CDG PAD_Inst_Cahe_writeData_data32 (.I(WIRE_Inst_Cahe_writeData_data[32]), .PAD(PO_Inst_Cahe_writeData_data[32]));
PDO02CDG PAD_Inst_Cahe_writeData_data33 (.I(WIRE_Inst_Cahe_writeData_data[33]), .PAD(PO_Inst_Cahe_writeData_data[33]));
PDO02CDG PAD_Inst_Cahe_writeData_data34 (.I(WIRE_Inst_Cahe_writeData_data[34]), .PAD(PO_Inst_Cahe_writeData_data[34]));
PDO02CDG PAD_Inst_Cahe_writeData_data35 (.I(WIRE_Inst_Cahe_writeData_data[35]), .PAD(PO_Inst_Cahe_writeData_data[35]));
PDO02CDG PAD_Inst_Cahe_writeData_data36 (.I(WIRE_Inst_Cahe_writeData_data[36]), .PAD(PO_Inst_Cahe_writeData_data[36]));
PDO02CDG PAD_Inst_Cahe_writeData_data37 (.I(WIRE_Inst_Cahe_writeData_data[37]), .PAD(PO_Inst_Cahe_writeData_data[37]));
PDO02CDG PAD_Inst_Cahe_writeData_data38 (.I(WIRE_Inst_Cahe_writeData_data[38]), .PAD(PO_Inst_Cahe_writeData_data[38]));
PDO02CDG PAD_Inst_Cahe_writeData_data39 (.I(WIRE_Inst_Cahe_writeData_data[39]), .PAD(PO_Inst_Cahe_writeData_data[39]));
PDO02CDG PAD_Inst_Cahe_writeData_data40 (.I(WIRE_Inst_Cahe_writeData_data[40]), .PAD(PO_Inst_Cahe_writeData_data[40]));
PDO02CDG PAD_Inst_Cahe_writeData_data41 (.I(WIRE_Inst_Cahe_writeData_data[41]), .PAD(PO_Inst_Cahe_writeData_data[41]));
PDO02CDG PAD_Inst_Cahe_writeData_data42 (.I(WIRE_Inst_Cahe_writeData_data[42]), .PAD(PO_Inst_Cahe_writeData_data[42]));
PDO02CDG PAD_Inst_Cahe_writeData_data43 (.I(WIRE_Inst_Cahe_writeData_data[43]), .PAD(PO_Inst_Cahe_writeData_data[43]));
PDO02CDG PAD_Inst_Cahe_writeData_data44 (.I(WIRE_Inst_Cahe_writeData_data[44]), .PAD(PO_Inst_Cahe_writeData_data[44]));
PDO02CDG PAD_Inst_Cahe_writeData_data45 (.I(WIRE_Inst_Cahe_writeData_data[45]), .PAD(PO_Inst_Cahe_writeData_data[45]));
PDO02CDG PAD_Inst_Cahe_writeData_data46 (.I(WIRE_Inst_Cahe_writeData_data[46]), .PAD(PO_Inst_Cahe_writeData_data[46]));
PDO02CDG PAD_Inst_Cahe_writeData_data47 (.I(WIRE_Inst_Cahe_writeData_data[47]), .PAD(PO_Inst_Cahe_writeData_data[47]));
PDO02CDG PAD_Inst_Cahe_writeData_data48 (.I(WIRE_Inst_Cahe_writeData_data[48]), .PAD(PO_Inst_Cahe_writeData_data[48]));
PDO02CDG PAD_Inst_Cahe_writeData_data49 (.I(WIRE_Inst_Cahe_writeData_data[49]), .PAD(PO_Inst_Cahe_writeData_data[49]));
PDO02CDG PAD_Inst_Cahe_writeData_data50 (.I(WIRE_Inst_Cahe_writeData_data[50]), .PAD(PO_Inst_Cahe_writeData_data[50]));
PDO02CDG PAD_Inst_Cahe_writeData_data51 (.I(WIRE_Inst_Cahe_writeData_data[51]), .PAD(PO_Inst_Cahe_writeData_data[51]));
PDO02CDG PAD_Inst_Cahe_writeData_data52 (.I(WIRE_Inst_Cahe_writeData_data[52]), .PAD(PO_Inst_Cahe_writeData_data[52]));
PDO02CDG PAD_Inst_Cahe_writeData_data53 (.I(WIRE_Inst_Cahe_writeData_data[53]), .PAD(PO_Inst_Cahe_writeData_data[53]));
PDO02CDG PAD_Inst_Cahe_writeData_data54 (.I(WIRE_Inst_Cahe_writeData_data[54]), .PAD(PO_Inst_Cahe_writeData_data[54]));
PDO02CDG PAD_Inst_Cahe_writeData_data55 (.I(WIRE_Inst_Cahe_writeData_data[55]), .PAD(PO_Inst_Cahe_writeData_data[55]));
PDO02CDG PAD_Inst_Cahe_writeData_data56 (.I(WIRE_Inst_Cahe_writeData_data[56]), .PAD(PO_Inst_Cahe_writeData_data[56]));
PDO02CDG PAD_Inst_Cahe_writeData_data57 (.I(WIRE_Inst_Cahe_writeData_data[57]), .PAD(PO_Inst_Cahe_writeData_data[57]));
PDO02CDG PAD_Inst_Cahe_writeData_data58 (.I(WIRE_Inst_Cahe_writeData_data[58]), .PAD(PO_Inst_Cahe_writeData_data[58]));
PDO02CDG PAD_Inst_Cahe_writeData_data59 (.I(WIRE_Inst_Cahe_writeData_data[59]), .PAD(PO_Inst_Cahe_writeData_data[59]));
PDO02CDG PAD_Inst_Cahe_writeData_data60 (.I(WIRE_Inst_Cahe_writeData_data[60]), .PAD(PO_Inst_Cahe_writeData_data[60]));
PDO02CDG PAD_Inst_Cahe_writeData_data61 (.I(WIRE_Inst_Cahe_writeData_data[61]), .PAD(PO_Inst_Cahe_writeData_data[61]));
PDO02CDG PAD_Inst_Cahe_writeData_data62 (.I(WIRE_Inst_Cahe_writeData_data[62]), .PAD(PO_Inst_Cahe_writeData_data[62]));
PDO02CDG PAD_Inst_Cahe_writeData_data63 (.I(WIRE_Inst_Cahe_writeData_data[63]), .PAD(PO_Inst_Cahe_writeData_data[63]));
PDO02CDG PAD_Inst_Cahe_writeData_data64 (.I(WIRE_Inst_Cahe_writeData_data[64]), .PAD(PO_Inst_Cahe_writeData_data[64]));
PDO02CDG PAD_Inst_Cahe_writeData_data65 (.I(WIRE_Inst_Cahe_writeData_data[65]), .PAD(PO_Inst_Cahe_writeData_data[65]));
PDO02CDG PAD_Inst_Cahe_writeData_data66 (.I(WIRE_Inst_Cahe_writeData_data[66]), .PAD(PO_Inst_Cahe_writeData_data[66]));
PDO02CDG PAD_Inst_Cahe_writeData_data67 (.I(WIRE_Inst_Cahe_writeData_data[67]), .PAD(PO_Inst_Cahe_writeData_data[67]));
PDO02CDG PAD_Inst_Cahe_writeData_data68 (.I(WIRE_Inst_Cahe_writeData_data[68]), .PAD(PO_Inst_Cahe_writeData_data[68]));
PDO02CDG PAD_Inst_Cahe_writeData_data69 (.I(WIRE_Inst_Cahe_writeData_data[69]), .PAD(PO_Inst_Cahe_writeData_data[69]));
PDO02CDG PAD_Inst_Cahe_writeData_data70 (.I(WIRE_Inst_Cahe_writeData_data[70]), .PAD(PO_Inst_Cahe_writeData_data[70]));
PDO02CDG PAD_Inst_Cahe_writeData_data71 (.I(WIRE_Inst_Cahe_writeData_data[71]), .PAD(PO_Inst_Cahe_writeData_data[71]));
PDO02CDG PAD_Inst_Cahe_writeData_data72 (.I(WIRE_Inst_Cahe_writeData_data[72]), .PAD(PO_Inst_Cahe_writeData_data[72]));
PDO02CDG PAD_Inst_Cahe_writeData_data73 (.I(WIRE_Inst_Cahe_writeData_data[73]), .PAD(PO_Inst_Cahe_writeData_data[73]));
PDO02CDG PAD_Inst_Cahe_writeData_data74 (.I(WIRE_Inst_Cahe_writeData_data[74]), .PAD(PO_Inst_Cahe_writeData_data[74]));
PDO02CDG PAD_Inst_Cahe_writeData_data75 (.I(WIRE_Inst_Cahe_writeData_data[75]), .PAD(PO_Inst_Cahe_writeData_data[75]));
PDO02CDG PAD_Inst_Cahe_writeData_data76 (.I(WIRE_Inst_Cahe_writeData_data[76]), .PAD(PO_Inst_Cahe_writeData_data[76]));
PDO02CDG PAD_Inst_Cahe_writeData_data77 (.I(WIRE_Inst_Cahe_writeData_data[77]), .PAD(PO_Inst_Cahe_writeData_data[77]));
PDO02CDG PAD_Inst_Cahe_writeData_data78 (.I(WIRE_Inst_Cahe_writeData_data[78]), .PAD(PO_Inst_Cahe_writeData_data[78]));
PDO02CDG PAD_Inst_Cahe_writeData_data79 (.I(WIRE_Inst_Cahe_writeData_data[79]), .PAD(PO_Inst_Cahe_writeData_data[79]));
PDO02CDG PAD_Inst_Cahe_writeData_data80 (.I(WIRE_Inst_Cahe_writeData_data[80]), .PAD(PO_Inst_Cahe_writeData_data[80]));
PDO02CDG PAD_Inst_Cahe_writeData_data81 (.I(WIRE_Inst_Cahe_writeData_data[81]), .PAD(PO_Inst_Cahe_writeData_data[81]));
PDO02CDG PAD_Inst_Cahe_writeData_data82 (.I(WIRE_Inst_Cahe_writeData_data[82]), .PAD(PO_Inst_Cahe_writeData_data[82]));
PDO02CDG PAD_Inst_Cahe_writeData_data83 (.I(WIRE_Inst_Cahe_writeData_data[83]), .PAD(PO_Inst_Cahe_writeData_data[83]));
PDO02CDG PAD_Inst_Cahe_writeData_data84 (.I(WIRE_Inst_Cahe_writeData_data[84]), .PAD(PO_Inst_Cahe_writeData_data[84]));
PDO02CDG PAD_Inst_Cahe_writeData_data85 (.I(WIRE_Inst_Cahe_writeData_data[85]), .PAD(PO_Inst_Cahe_writeData_data[85]));
PDO02CDG PAD_Inst_Cahe_writeData_data86 (.I(WIRE_Inst_Cahe_writeData_data[86]), .PAD(PO_Inst_Cahe_writeData_data[86]));
PDO02CDG PAD_Inst_Cahe_writeData_data87 (.I(WIRE_Inst_Cahe_writeData_data[87]), .PAD(PO_Inst_Cahe_writeData_data[87]));
PDO02CDG PAD_Inst_Cahe_writeData_data88 (.I(WIRE_Inst_Cahe_writeData_data[88]), .PAD(PO_Inst_Cahe_writeData_data[88]));
PDO02CDG PAD_Inst_Cahe_writeData_data89 (.I(WIRE_Inst_Cahe_writeData_data[89]), .PAD(PO_Inst_Cahe_writeData_data[89]));
PDO02CDG PAD_Inst_Cahe_writeData_data90 (.I(WIRE_Inst_Cahe_writeData_data[90]), .PAD(PO_Inst_Cahe_writeData_data[90]));
PDO02CDG PAD_Inst_Cahe_writeData_data91 (.I(WIRE_Inst_Cahe_writeData_data[91]), .PAD(PO_Inst_Cahe_writeData_data[91]));
PDO02CDG PAD_Inst_Cahe_writeData_data92 (.I(WIRE_Inst_Cahe_writeData_data[92]), .PAD(PO_Inst_Cahe_writeData_data[92]));
PDO02CDG PAD_Inst_Cahe_writeData_data93 (.I(WIRE_Inst_Cahe_writeData_data[93]), .PAD(PO_Inst_Cahe_writeData_data[93]));
PDO02CDG PAD_Inst_Cahe_writeData_data94 (.I(WIRE_Inst_Cahe_writeData_data[94]), .PAD(PO_Inst_Cahe_writeData_data[94]));
PDO02CDG PAD_Inst_Cahe_writeData_data95 (.I(WIRE_Inst_Cahe_writeData_data[95]), .PAD(PO_Inst_Cahe_writeData_data[95]));
PDO02CDG PAD_Inst_Cahe_writeData_data96 (.I(WIRE_Inst_Cahe_writeData_data[96]), .PAD(PO_Inst_Cahe_writeData_data[96]));
PDO02CDG PAD_Inst_Cahe_writeData_data97 (.I(WIRE_Inst_Cahe_writeData_data[97]), .PAD(PO_Inst_Cahe_writeData_data[97]));
PDO02CDG PAD_Inst_Cahe_writeData_data98 (.I(WIRE_Inst_Cahe_writeData_data[98]), .PAD(PO_Inst_Cahe_writeData_data[98]));
PDO02CDG PAD_Inst_Cahe_writeData_data99 (.I(WIRE_Inst_Cahe_writeData_data[99]), .PAD(PO_Inst_Cahe_writeData_data[99]));
PDO02CDG PAD_Inst_Cahe_writeData_data100 (.I(WIRE_Inst_Cahe_writeData_data[100]), .PAD(PO_Inst_Cahe_writeData_data[100]));
PDO02CDG PAD_Inst_Cahe_writeData_data101 (.I(WIRE_Inst_Cahe_writeData_data[101]), .PAD(PO_Inst_Cahe_writeData_data[101]));
PDO02CDG PAD_Inst_Cahe_writeData_data102 (.I(WIRE_Inst_Cahe_writeData_data[102]), .PAD(PO_Inst_Cahe_writeData_data[102]));
PDO02CDG PAD_Inst_Cahe_writeData_data103 (.I(WIRE_Inst_Cahe_writeData_data[103]), .PAD(PO_Inst_Cahe_writeData_data[103]));
PDO02CDG PAD_Inst_Cahe_writeData_data104 (.I(WIRE_Inst_Cahe_writeData_data[104]), .PAD(PO_Inst_Cahe_writeData_data[104]));
PDO02CDG PAD_Inst_Cahe_writeData_data105 (.I(WIRE_Inst_Cahe_writeData_data[105]), .PAD(PO_Inst_Cahe_writeData_data[105]));
PDO02CDG PAD_Inst_Cahe_writeData_data106 (.I(WIRE_Inst_Cahe_writeData_data[106]), .PAD(PO_Inst_Cahe_writeData_data[106]));
PDO02CDG PAD_Inst_Cahe_writeData_data107 (.I(WIRE_Inst_Cahe_writeData_data[107]), .PAD(PO_Inst_Cahe_writeData_data[107]));
PDO02CDG PAD_Inst_Cahe_writeData_data108 (.I(WIRE_Inst_Cahe_writeData_data[108]), .PAD(PO_Inst_Cahe_writeData_data[108]));
PDO02CDG PAD_Inst_Cahe_writeData_data109 (.I(WIRE_Inst_Cahe_writeData_data[109]), .PAD(PO_Inst_Cahe_writeData_data[109]));
PDO02CDG PAD_Inst_Cahe_writeData_data110 (.I(WIRE_Inst_Cahe_writeData_data[110]), .PAD(PO_Inst_Cahe_writeData_data[110]));
PDO02CDG PAD_Inst_Cahe_writeData_data111 (.I(WIRE_Inst_Cahe_writeData_data[111]), .PAD(PO_Inst_Cahe_writeData_data[111]));
PDO02CDG PAD_Inst_Cahe_writeData_data112 (.I(WIRE_Inst_Cahe_writeData_data[112]), .PAD(PO_Inst_Cahe_writeData_data[112]));
PDO02CDG PAD_Inst_Cahe_writeData_data113 (.I(WIRE_Inst_Cahe_writeData_data[113]), .PAD(PO_Inst_Cahe_writeData_data[113]));
PDO02CDG PAD_Inst_Cahe_writeData_data114 (.I(WIRE_Inst_Cahe_writeData_data[114]), .PAD(PO_Inst_Cahe_writeData_data[114]));
PDO02CDG PAD_Inst_Cahe_writeData_data115 (.I(WIRE_Inst_Cahe_writeData_data[115]), .PAD(PO_Inst_Cahe_writeData_data[115]));
PDO02CDG PAD_Inst_Cahe_writeData_data116 (.I(WIRE_Inst_Cahe_writeData_data[116]), .PAD(PO_Inst_Cahe_writeData_data[116]));
PDO02CDG PAD_Inst_Cahe_writeData_data117 (.I(WIRE_Inst_Cahe_writeData_data[117]), .PAD(PO_Inst_Cahe_writeData_data[117]));
PDO02CDG PAD_Inst_Cahe_writeData_data118 (.I(WIRE_Inst_Cahe_writeData_data[118]), .PAD(PO_Inst_Cahe_writeData_data[118]));
PDO02CDG PAD_Inst_Cahe_writeData_data119 (.I(WIRE_Inst_Cahe_writeData_data[119]), .PAD(PO_Inst_Cahe_writeData_data[119]));
PDO02CDG PAD_Inst_Cahe_writeData_data120 (.I(WIRE_Inst_Cahe_writeData_data[120]), .PAD(PO_Inst_Cahe_writeData_data[120]));
PDO02CDG PAD_Inst_Cahe_writeData_data121 (.I(WIRE_Inst_Cahe_writeData_data[121]), .PAD(PO_Inst_Cahe_writeData_data[121]));
PDO02CDG PAD_Inst_Cahe_writeData_data122 (.I(WIRE_Inst_Cahe_writeData_data[122]), .PAD(PO_Inst_Cahe_writeData_data[122]));
PDO02CDG PAD_Inst_Cahe_writeData_data123 (.I(WIRE_Inst_Cahe_writeData_data[123]), .PAD(PO_Inst_Cahe_writeData_data[123]));
PDO02CDG PAD_Inst_Cahe_writeData_data124 (.I(WIRE_Inst_Cahe_writeData_data[124]), .PAD(PO_Inst_Cahe_writeData_data[124]));
PDO02CDG PAD_Inst_Cahe_writeData_data125 (.I(WIRE_Inst_Cahe_writeData_data[125]), .PAD(PO_Inst_Cahe_writeData_data[125]));
PDO02CDG PAD_Inst_Cahe_writeData_data126 (.I(WIRE_Inst_Cahe_writeData_data[126]), .PAD(PO_Inst_Cahe_writeData_data[126]));
PDO02CDG PAD_Inst_Cahe_writeData_data127 (.I(WIRE_Inst_Cahe_writeData_data[127]), .PAD(PO_Inst_Cahe_writeData_data[127]));

PDO02CDG PAD_Inst_Cahe_writeData_strb0 (.I(WIRE_Inst_Cahe_writeData_strb[0]), .PAD(PO_Inst_Cahe_writeData_strb[0]));
PDO02CDG PAD_Inst_Cahe_writeData_strb1 (.I(WIRE_Inst_Cahe_writeData_strb[1]), .PAD(PO_Inst_Cahe_writeData_strb[1]));
PDO02CDG PAD_Inst_Cahe_writeData_strb2 (.I(WIRE_Inst_Cahe_writeData_strb[2]), .PAD(PO_Inst_Cahe_writeData_strb[2]));
PDO02CDG PAD_Inst_Cahe_writeData_strb3 (.I(WIRE_Inst_Cahe_writeData_strb[3]), .PAD(PO_Inst_Cahe_writeData_strb[3]));
PDO02CDG PAD_Inst_Cahe_writeData_strb4 (.I(WIRE_Inst_Cahe_writeData_strb[4]), .PAD(PO_Inst_Cahe_writeData_strb[4]));
PDO02CDG PAD_Inst_Cahe_writeData_strb5 (.I(WIRE_Inst_Cahe_writeData_strb[5]), .PAD(PO_Inst_Cahe_writeData_strb[5]));
PDO02CDG PAD_Inst_Cahe_writeData_strb6 (.I(WIRE_Inst_Cahe_writeData_strb[6]), .PAD(PO_Inst_Cahe_writeData_strb[6]));
PDO02CDG PAD_Inst_Cahe_writeData_strb7 (.I(WIRE_Inst_Cahe_writeData_strb[7]), .PAD(PO_Inst_Cahe_writeData_strb[7]));
PDO02CDG PAD_Inst_Cahe_writeData_strb8 (.I(WIRE_Inst_Cahe_writeData_strb[8]), .PAD(PO_Inst_Cahe_writeData_strb[8]));
PDO02CDG PAD_Inst_Cahe_writeData_strb9 (.I(WIRE_Inst_Cahe_writeData_strb[9]), .PAD(PO_Inst_Cahe_writeData_strb[9]));
PDO02CDG PAD_Inst_Cahe_writeData_strb10 (.I(WIRE_Inst_Cahe_writeData_strb[10]), .PAD(PO_Inst_Cahe_writeData_strb[10]));
PDO02CDG PAD_Inst_Cahe_writeData_strb11 (.I(WIRE_Inst_Cahe_writeData_strb[11]), .PAD(PO_Inst_Cahe_writeData_strb[11]));
PDO02CDG PAD_Inst_Cahe_writeData_strb12 (.I(WIRE_Inst_Cahe_writeData_strb[12]), .PAD(PO_Inst_Cahe_writeData_strb[12]));
PDO02CDG PAD_Inst_Cahe_writeData_strb13 (.I(WIRE_Inst_Cahe_writeData_strb[13]), .PAD(PO_Inst_Cahe_writeData_strb[13]));
PDO02CDG PAD_Inst_Cahe_writeData_strb14 (.I(WIRE_Inst_Cahe_writeData_strb[14]), .PAD(PO_Inst_Cahe_writeData_strb[14]));
PDO02CDG PAD_Inst_Cahe_writeData_strb15 (.I(WIRE_Inst_Cahe_writeData_strb[15]), .PAD(PO_Inst_Cahe_writeData_strb[15]));

PDO02CDG PAD_Inst_Cahe_writeData_valid (.I(WIRE_Inst_Cahe_writeData_valid), .PAD(PO_Inst_Cahe_writeData_valid));
PDO02CDG PAD_Inst_Cahe_writeResp_ready (.I(WIRE_Inst_Cahe_writeResp_ready), .PAD(PO_Inst_Cahe_writeResp_ready));

// CORNER3

PDO02CDG PAD_Data_Cahe_readAddr_addr0 (.I(WIRE_Data_Cahe_readAddr_addr[0]), .PAD(PO_Data_Cahe_readAddr_addr[0]));
PDO02CDG PAD_Data_Cahe_readAddr_addr1 (.I(WIRE_Data_Cahe_readAddr_addr[1]), .PAD(PO_Data_Cahe_readAddr_addr[1]));
PDO02CDG PAD_Data_Cahe_readAddr_addr2 (.I(WIRE_Data_Cahe_readAddr_addr[2]), .PAD(PO_Data_Cahe_readAddr_addr[2]));
PDO02CDG PAD_Data_Cahe_readAddr_addr3 (.I(WIRE_Data_Cahe_readAddr_addr[3]), .PAD(PO_Data_Cahe_readAddr_addr[3]));
PDO02CDG PAD_Data_Cahe_readAddr_addr4 (.I(WIRE_Data_Cahe_readAddr_addr[4]), .PAD(PO_Data_Cahe_readAddr_addr[4]));
PDO02CDG PAD_Data_Cahe_readAddr_addr5 (.I(WIRE_Data_Cahe_readAddr_addr[5]), .PAD(PO_Data_Cahe_readAddr_addr[5]));
PDO02CDG PAD_Data_Cahe_readAddr_addr6 (.I(WIRE_Data_Cahe_readAddr_addr[6]), .PAD(PO_Data_Cahe_readAddr_addr[6]));
PDO02CDG PAD_Data_Cahe_readAddr_addr7 (.I(WIRE_Data_Cahe_readAddr_addr[7]), .PAD(PO_Data_Cahe_readAddr_addr[7]));
PDO02CDG PAD_Data_Cahe_readAddr_addr8 (.I(WIRE_Data_Cahe_readAddr_addr[8]), .PAD(PO_Data_Cahe_readAddr_addr[8]));
PDO02CDG PAD_Data_Cahe_readAddr_addr9 (.I(WIRE_Data_Cahe_readAddr_addr[9]), .PAD(PO_Data_Cahe_readAddr_addr[9]));
PDO02CDG PAD_Data_Cahe_readAddr_addr10 (.I(WIRE_Data_Cahe_readAddr_addr[10]), .PAD(PO_Data_Cahe_readAddr_addr[10]));
PDO02CDG PAD_Data_Cahe_readAddr_addr11 (.I(WIRE_Data_Cahe_readAddr_addr[11]), .PAD(PO_Data_Cahe_readAddr_addr[11]));
PDO02CDG PAD_Data_Cahe_readAddr_addr12 (.I(WIRE_Data_Cahe_readAddr_addr[12]), .PAD(PO_Data_Cahe_readAddr_addr[12]));
PDO02CDG PAD_Data_Cahe_readAddr_addr13 (.I(WIRE_Data_Cahe_readAddr_addr[13]), .PAD(PO_Data_Cahe_readAddr_addr[13]));
PDO02CDG PAD_Data_Cahe_readAddr_addr14 (.I(WIRE_Data_Cahe_readAddr_addr[14]), .PAD(PO_Data_Cahe_readAddr_addr[14]));
PDO02CDG PAD_Data_Cahe_readAddr_addr15 (.I(WIRE_Data_Cahe_readAddr_addr[15]), .PAD(PO_Data_Cahe_readAddr_addr[15]));
PDO02CDG PAD_Data_Cahe_readAddr_addr16 (.I(WIRE_Data_Cahe_readAddr_addr[16]), .PAD(PO_Data_Cahe_readAddr_addr[16]));
PDO02CDG PAD_Data_Cahe_readAddr_addr17 (.I(WIRE_Data_Cahe_readAddr_addr[17]), .PAD(PO_Data_Cahe_readAddr_addr[17]));
PDO02CDG PAD_Data_Cahe_readAddr_addr18 (.I(WIRE_Data_Cahe_readAddr_addr[18]), .PAD(PO_Data_Cahe_readAddr_addr[18]));
PDO02CDG PAD_Data_Cahe_readAddr_addr19 (.I(WIRE_Data_Cahe_readAddr_addr[19]), .PAD(PO_Data_Cahe_readAddr_addr[19]));
PDO02CDG PAD_Data_Cahe_readAddr_addr20 (.I(WIRE_Data_Cahe_readAddr_addr[20]), .PAD(PO_Data_Cahe_readAddr_addr[20]));
PDO02CDG PAD_Data_Cahe_readAddr_addr21 (.I(WIRE_Data_Cahe_readAddr_addr[21]), .PAD(PO_Data_Cahe_readAddr_addr[21]));
PDO02CDG PAD_Data_Cahe_readAddr_addr22 (.I(WIRE_Data_Cahe_readAddr_addr[22]), .PAD(PO_Data_Cahe_readAddr_addr[22]));
PDO02CDG PAD_Data_Cahe_readAddr_addr23 (.I(WIRE_Data_Cahe_readAddr_addr[23]), .PAD(PO_Data_Cahe_readAddr_addr[23]));
PDO02CDG PAD_Data_Cahe_readAddr_addr24 (.I(WIRE_Data_Cahe_readAddr_addr[24]), .PAD(PO_Data_Cahe_readAddr_addr[24]));
PDO02CDG PAD_Data_Cahe_readAddr_addr25 (.I(WIRE_Data_Cahe_readAddr_addr[25]), .PAD(PO_Data_Cahe_readAddr_addr[25]));
PDO02CDG PAD_Data_Cahe_readAddr_addr26 (.I(WIRE_Data_Cahe_readAddr_addr[26]), .PAD(PO_Data_Cahe_readAddr_addr[26]));
PDO02CDG PAD_Data_Cahe_readAddr_addr27 (.I(WIRE_Data_Cahe_readAddr_addr[27]), .PAD(PO_Data_Cahe_readAddr_addr[27]));
PDO02CDG PAD_Data_Cahe_readAddr_addr28 (.I(WIRE_Data_Cahe_readAddr_addr[28]), .PAD(PO_Data_Cahe_readAddr_addr[28]));
PDO02CDG PAD_Data_Cahe_readAddr_addr29 (.I(WIRE_Data_Cahe_readAddr_addr[29]), .PAD(PO_Data_Cahe_readAddr_addr[29]));
PDO02CDG PAD_Data_Cahe_readAddr_addr30 (.I(WIRE_Data_Cahe_readAddr_addr[30]), .PAD(PO_Data_Cahe_readAddr_addr[30]));
PDO02CDG PAD_Data_Cahe_readAddr_addr31 (.I(WIRE_Data_Cahe_readAddr_addr[31]), .PAD(PO_Data_Cahe_readAddr_addr[31]));

PDO02CDG PAD_Data_Cahe_readAddr_valid  (.I(WIRE_Data_Cahe_readAddr_valid), .PAD(PO_Data_Cahe_readAddr_valid));
PDO02CDG PAD_Data_Cahe_readData_ready  (.I(WIRE_Data_Cahe_readData_ready), .PAD(PO_Data_Cahe_readData_ready));

PDO02CDG PAD_Data_Cahe_writeAddr_addr0 (.I(WIRE_Data_Cahe_writeAddr_addr[0]), .PAD(PO_Data_Cahe_writeAddr_addr[0]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr1 (.I(WIRE_Data_Cahe_writeAddr_addr[1]), .PAD(PO_Data_Cahe_writeAddr_addr[1]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr2 (.I(WIRE_Data_Cahe_writeAddr_addr[2]), .PAD(PO_Data_Cahe_writeAddr_addr[2]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr3 (.I(WIRE_Data_Cahe_writeAddr_addr[3]), .PAD(PO_Data_Cahe_writeAddr_addr[3]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr4 (.I(WIRE_Data_Cahe_writeAddr_addr[4]), .PAD(PO_Data_Cahe_writeAddr_addr[4]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr5 (.I(WIRE_Data_Cahe_writeAddr_addr[5]), .PAD(PO_Data_Cahe_writeAddr_addr[5]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr6 (.I(WIRE_Data_Cahe_writeAddr_addr[6]), .PAD(PO_Data_Cahe_writeAddr_addr[6]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr7 (.I(WIRE_Data_Cahe_writeAddr_addr[7]), .PAD(PO_Data_Cahe_writeAddr_addr[7]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr8 (.I(WIRE_Data_Cahe_writeAddr_addr[8]), .PAD(PO_Data_Cahe_writeAddr_addr[8]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr9 (.I(WIRE_Data_Cahe_writeAddr_addr[9]), .PAD(PO_Data_Cahe_writeAddr_addr[9]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr10 (.I(WIRE_Data_Cahe_writeAddr_addr[10]), .PAD(PO_Data_Cahe_writeAddr_addr[10]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr11 (.I(WIRE_Data_Cahe_writeAddr_addr[11]), .PAD(PO_Data_Cahe_writeAddr_addr[11]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr12 (.I(WIRE_Data_Cahe_writeAddr_addr[12]), .PAD(PO_Data_Cahe_writeAddr_addr[12]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr13 (.I(WIRE_Data_Cahe_writeAddr_addr[13]), .PAD(PO_Data_Cahe_writeAddr_addr[13]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr14 (.I(WIRE_Data_Cahe_writeAddr_addr[14]), .PAD(PO_Data_Cahe_writeAddr_addr[14]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr15 (.I(WIRE_Data_Cahe_writeAddr_addr[15]), .PAD(PO_Data_Cahe_writeAddr_addr[15]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr16 (.I(WIRE_Data_Cahe_writeAddr_addr[16]), .PAD(PO_Data_Cahe_writeAddr_addr[16]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr17 (.I(WIRE_Data_Cahe_writeAddr_addr[17]), .PAD(PO_Data_Cahe_writeAddr_addr[17]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr18 (.I(WIRE_Data_Cahe_writeAddr_addr[18]), .PAD(PO_Data_Cahe_writeAddr_addr[18]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr19 (.I(WIRE_Data_Cahe_writeAddr_addr[19]), .PAD(PO_Data_Cahe_writeAddr_addr[19]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr20 (.I(WIRE_Data_Cahe_writeAddr_addr[20]), .PAD(PO_Data_Cahe_writeAddr_addr[20]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr21 (.I(WIRE_Data_Cahe_writeAddr_addr[21]), .PAD(PO_Data_Cahe_writeAddr_addr[21]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr22 (.I(WIRE_Data_Cahe_writeAddr_addr[22]), .PAD(PO_Data_Cahe_writeAddr_addr[22]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr23 (.I(WIRE_Data_Cahe_writeAddr_addr[23]), .PAD(PO_Data_Cahe_writeAddr_addr[23]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr24 (.I(WIRE_Data_Cahe_writeAddr_addr[24]), .PAD(PO_Data_Cahe_writeAddr_addr[24]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr25 (.I(WIRE_Data_Cahe_writeAddr_addr[25]), .PAD(PO_Data_Cahe_writeAddr_addr[25]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr26 (.I(WIRE_Data_Cahe_writeAddr_addr[26]), .PAD(PO_Data_Cahe_writeAddr_addr[26]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr27 (.I(WIRE_Data_Cahe_writeAddr_addr[27]), .PAD(PO_Data_Cahe_writeAddr_addr[27]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr28 (.I(WIRE_Data_Cahe_writeAddr_addr[28]), .PAD(PO_Data_Cahe_writeAddr_addr[28]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr29 (.I(WIRE_Data_Cahe_writeAddr_addr[29]), .PAD(PO_Data_Cahe_writeAddr_addr[29]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr30 (.I(WIRE_Data_Cahe_writeAddr_addr[30]), .PAD(PO_Data_Cahe_writeAddr_addr[30]));
PDO02CDG PAD_Data_Cahe_writeAddr_addr31 (.I(WIRE_Data_Cahe_writeAddr_addr[31]), .PAD(PO_Data_Cahe_writeAddr_addr[31]));

PDO02CDG PAD_Data_Cahe_writeAddr_valid (.I(WIRE_Data_Cahe_writeAddr_valid), .PAD(PO_Data_Cahe_writeAddr_valid));

PDO02CDG PAD_Data_Cahe_writeData_data0 (.I(WIRE_Data_Cahe_writeData_data[0]), .PAD(PO_Data_Cahe_writeData_data[0]));
PDO02CDG PAD_Data_Cahe_writeData_data1 (.I(WIRE_Data_Cahe_writeData_data[1]), .PAD(PO_Data_Cahe_writeData_data[1]));
PDO02CDG PAD_Data_Cahe_writeData_data2 (.I(WIRE_Data_Cahe_writeData_data[2]), .PAD(PO_Data_Cahe_writeData_data[2]));
PDO02CDG PAD_Data_Cahe_writeData_data3 (.I(WIRE_Data_Cahe_writeData_data[3]), .PAD(PO_Data_Cahe_writeData_data[3]));
PDO02CDG PAD_Data_Cahe_writeData_data4 (.I(WIRE_Data_Cahe_writeData_data[4]), .PAD(PO_Data_Cahe_writeData_data[4]));
PDO02CDG PAD_Data_Cahe_writeData_data5 (.I(WIRE_Data_Cahe_writeData_data[5]), .PAD(PO_Data_Cahe_writeData_data[5]));
PDO02CDG PAD_Data_Cahe_writeData_data6 (.I(WIRE_Data_Cahe_writeData_data[6]), .PAD(PO_Data_Cahe_writeData_data[6]));
PDO02CDG PAD_Data_Cahe_writeData_data7 (.I(WIRE_Data_Cahe_writeData_data[7]), .PAD(PO_Data_Cahe_writeData_data[7]));
PDO02CDG PAD_Data_Cahe_writeData_data8 (.I(WIRE_Data_Cahe_writeData_data[8]), .PAD(PO_Data_Cahe_writeData_data[8]));
PDO02CDG PAD_Data_Cahe_writeData_data9 (.I(WIRE_Data_Cahe_writeData_data[9]), .PAD(PO_Data_Cahe_writeData_data[9]));
PDO02CDG PAD_Data_Cahe_writeData_data10 (.I(WIRE_Data_Cahe_writeData_data[10]), .PAD(PO_Data_Cahe_writeData_data[10]));
PDO02CDG PAD_Data_Cahe_writeData_data11 (.I(WIRE_Data_Cahe_writeData_data[11]), .PAD(PO_Data_Cahe_writeData_data[11]));
PDO02CDG PAD_Data_Cahe_writeData_data12 (.I(WIRE_Data_Cahe_writeData_data[12]), .PAD(PO_Data_Cahe_writeData_data[12]));
PDO02CDG PAD_Data_Cahe_writeData_data13 (.I(WIRE_Data_Cahe_writeData_data[13]), .PAD(PO_Data_Cahe_writeData_data[13]));
PDO02CDG PAD_Data_Cahe_writeData_data14 (.I(WIRE_Data_Cahe_writeData_data[14]), .PAD(PO_Data_Cahe_writeData_data[14]));
PDO02CDG PAD_Data_Cahe_writeData_data15 (.I(WIRE_Data_Cahe_writeData_data[15]), .PAD(PO_Data_Cahe_writeData_data[15]));
PDO02CDG PAD_Data_Cahe_writeData_data16 (.I(WIRE_Data_Cahe_writeData_data[16]), .PAD(PO_Data_Cahe_writeData_data[16]));
PDO02CDG PAD_Data_Cahe_writeData_data17 (.I(WIRE_Data_Cahe_writeData_data[17]), .PAD(PO_Data_Cahe_writeData_data[17]));
PDO02CDG PAD_Data_Cahe_writeData_data18 (.I(WIRE_Data_Cahe_writeData_data[18]), .PAD(PO_Data_Cahe_writeData_data[18]));
PDO02CDG PAD_Data_Cahe_writeData_data19 (.I(WIRE_Data_Cahe_writeData_data[19]), .PAD(PO_Data_Cahe_writeData_data[19]));
PDO02CDG PAD_Data_Cahe_writeData_data20 (.I(WIRE_Data_Cahe_writeData_data[20]), .PAD(PO_Data_Cahe_writeData_data[20]));
PDO02CDG PAD_Data_Cahe_writeData_data21 (.I(WIRE_Data_Cahe_writeData_data[21]), .PAD(PO_Data_Cahe_writeData_data[21]));
PDO02CDG PAD_Data_Cahe_writeData_data22 (.I(WIRE_Data_Cahe_writeData_data[22]), .PAD(PO_Data_Cahe_writeData_data[22]));
PDO02CDG PAD_Data_Cahe_writeData_data23 (.I(WIRE_Data_Cahe_writeData_data[23]), .PAD(PO_Data_Cahe_writeData_data[23]));
PDO02CDG PAD_Data_Cahe_writeData_data24 (.I(WIRE_Data_Cahe_writeData_data[24]), .PAD(PO_Data_Cahe_writeData_data[24]));
PDO02CDG PAD_Data_Cahe_writeData_data25 (.I(WIRE_Data_Cahe_writeData_data[25]), .PAD(PO_Data_Cahe_writeData_data[25]));
PDO02CDG PAD_Data_Cahe_writeData_data26 (.I(WIRE_Data_Cahe_writeData_data[26]), .PAD(PO_Data_Cahe_writeData_data[26]));
PDO02CDG PAD_Data_Cahe_writeData_data27 (.I(WIRE_Data_Cahe_writeData_data[27]), .PAD(PO_Data_Cahe_writeData_data[27]));
PDO02CDG PAD_Data_Cahe_writeData_data28 (.I(WIRE_Data_Cahe_writeData_data[28]), .PAD(PO_Data_Cahe_writeData_data[28]));
PDO02CDG PAD_Data_Cahe_writeData_data29 (.I(WIRE_Data_Cahe_writeData_data[29]), .PAD(PO_Data_Cahe_writeData_data[29]));
PDO02CDG PAD_Data_Cahe_writeData_data30 (.I(WIRE_Data_Cahe_writeData_data[30]), .PAD(PO_Data_Cahe_writeData_data[30]));
PDO02CDG PAD_Data_Cahe_writeData_data31 (.I(WIRE_Data_Cahe_writeData_data[31]), .PAD(PO_Data_Cahe_writeData_data[31]));
PDO02CDG PAD_Data_Cahe_writeData_data32 (.I(WIRE_Data_Cahe_writeData_data[32]), .PAD(PO_Data_Cahe_writeData_data[32]));
PDO02CDG PAD_Data_Cahe_writeData_data33 (.I(WIRE_Data_Cahe_writeData_data[33]), .PAD(PO_Data_Cahe_writeData_data[33]));
PDO02CDG PAD_Data_Cahe_writeData_data34 (.I(WIRE_Data_Cahe_writeData_data[34]), .PAD(PO_Data_Cahe_writeData_data[34]));
PDO02CDG PAD_Data_Cahe_writeData_data35 (.I(WIRE_Data_Cahe_writeData_data[35]), .PAD(PO_Data_Cahe_writeData_data[35]));
PDO02CDG PAD_Data_Cahe_writeData_data36 (.I(WIRE_Data_Cahe_writeData_data[36]), .PAD(PO_Data_Cahe_writeData_data[36]));
PDO02CDG PAD_Data_Cahe_writeData_data37 (.I(WIRE_Data_Cahe_writeData_data[37]), .PAD(PO_Data_Cahe_writeData_data[37]));
PDO02CDG PAD_Data_Cahe_writeData_data38 (.I(WIRE_Data_Cahe_writeData_data[38]), .PAD(PO_Data_Cahe_writeData_data[38]));
PDO02CDG PAD_Data_Cahe_writeData_data39 (.I(WIRE_Data_Cahe_writeData_data[39]), .PAD(PO_Data_Cahe_writeData_data[39]));
PDO02CDG PAD_Data_Cahe_writeData_data40 (.I(WIRE_Data_Cahe_writeData_data[40]), .PAD(PO_Data_Cahe_writeData_data[40]));
PDO02CDG PAD_Data_Cahe_writeData_data41 (.I(WIRE_Data_Cahe_writeData_data[41]), .PAD(PO_Data_Cahe_writeData_data[41]));
PDO02CDG PAD_Data_Cahe_writeData_data42 (.I(WIRE_Data_Cahe_writeData_data[42]), .PAD(PO_Data_Cahe_writeData_data[42]));
PDO02CDG PAD_Data_Cahe_writeData_data43 (.I(WIRE_Data_Cahe_writeData_data[43]), .PAD(PO_Data_Cahe_writeData_data[43]));
PDO02CDG PAD_Data_Cahe_writeData_data44 (.I(WIRE_Data_Cahe_writeData_data[44]), .PAD(PO_Data_Cahe_writeData_data[44]));
PDO02CDG PAD_Data_Cahe_writeData_data45 (.I(WIRE_Data_Cahe_writeData_data[45]), .PAD(PO_Data_Cahe_writeData_data[45]));
PDO02CDG PAD_Data_Cahe_writeData_data46 (.I(WIRE_Data_Cahe_writeData_data[46]), .PAD(PO_Data_Cahe_writeData_data[46]));
PDO02CDG PAD_Data_Cahe_writeData_data47 (.I(WIRE_Data_Cahe_writeData_data[47]), .PAD(PO_Data_Cahe_writeData_data[47]));
PDO02CDG PAD_Data_Cahe_writeData_data48 (.I(WIRE_Data_Cahe_writeData_data[48]), .PAD(PO_Data_Cahe_writeData_data[48]));
PDO02CDG PAD_Data_Cahe_writeData_data49 (.I(WIRE_Data_Cahe_writeData_data[49]), .PAD(PO_Data_Cahe_writeData_data[49]));
PDO02CDG PAD_Data_Cahe_writeData_data50 (.I(WIRE_Data_Cahe_writeData_data[50]), .PAD(PO_Data_Cahe_writeData_data[50]));
PDO02CDG PAD_Data_Cahe_writeData_data51 (.I(WIRE_Data_Cahe_writeData_data[51]), .PAD(PO_Data_Cahe_writeData_data[51]));
PDO02CDG PAD_Data_Cahe_writeData_data52 (.I(WIRE_Data_Cahe_writeData_data[52]), .PAD(PO_Data_Cahe_writeData_data[52]));
PDO02CDG PAD_Data_Cahe_writeData_data53 (.I(WIRE_Data_Cahe_writeData_data[53]), .PAD(PO_Data_Cahe_writeData_data[53]));
PDO02CDG PAD_Data_Cahe_writeData_data54 (.I(WIRE_Data_Cahe_writeData_data[54]), .PAD(PO_Data_Cahe_writeData_data[54]));
PDO02CDG PAD_Data_Cahe_writeData_data55 (.I(WIRE_Data_Cahe_writeData_data[55]), .PAD(PO_Data_Cahe_writeData_data[55]));
PDO02CDG PAD_Data_Cahe_writeData_data56 (.I(WIRE_Data_Cahe_writeData_data[56]), .PAD(PO_Data_Cahe_writeData_data[56]));
PDO02CDG PAD_Data_Cahe_writeData_data57 (.I(WIRE_Data_Cahe_writeData_data[57]), .PAD(PO_Data_Cahe_writeData_data[57]));
PDO02CDG PAD_Data_Cahe_writeData_data58 (.I(WIRE_Data_Cahe_writeData_data[58]), .PAD(PO_Data_Cahe_writeData_data[58]));
PDO02CDG PAD_Data_Cahe_writeData_data59 (.I(WIRE_Data_Cahe_writeData_data[59]), .PAD(PO_Data_Cahe_writeData_data[59]));
PDO02CDG PAD_Data_Cahe_writeData_data60 (.I(WIRE_Data_Cahe_writeData_data[60]), .PAD(PO_Data_Cahe_writeData_data[60]));
PDO02CDG PAD_Data_Cahe_writeData_data61 (.I(WIRE_Data_Cahe_writeData_data[61]), .PAD(PO_Data_Cahe_writeData_data[61]));
PDO02CDG PAD_Data_Cahe_writeData_data62 (.I(WIRE_Data_Cahe_writeData_data[62]), .PAD(PO_Data_Cahe_writeData_data[62]));
PDO02CDG PAD_Data_Cahe_writeData_data63 (.I(WIRE_Data_Cahe_writeData_data[63]), .PAD(PO_Data_Cahe_writeData_data[63]));
PDO02CDG PAD_Data_Cahe_writeData_data64 (.I(WIRE_Data_Cahe_writeData_data[64]), .PAD(PO_Data_Cahe_writeData_data[64]));
PDO02CDG PAD_Data_Cahe_writeData_data65 (.I(WIRE_Data_Cahe_writeData_data[65]), .PAD(PO_Data_Cahe_writeData_data[65]));
PDO02CDG PAD_Data_Cahe_writeData_data66 (.I(WIRE_Data_Cahe_writeData_data[66]), .PAD(PO_Data_Cahe_writeData_data[66]));
PDO02CDG PAD_Data_Cahe_writeData_data67 (.I(WIRE_Data_Cahe_writeData_data[67]), .PAD(PO_Data_Cahe_writeData_data[67]));
PDO02CDG PAD_Data_Cahe_writeData_data68 (.I(WIRE_Data_Cahe_writeData_data[68]), .PAD(PO_Data_Cahe_writeData_data[68]));
PDO02CDG PAD_Data_Cahe_writeData_data69 (.I(WIRE_Data_Cahe_writeData_data[69]), .PAD(PO_Data_Cahe_writeData_data[69]));
PDO02CDG PAD_Data_Cahe_writeData_data70 (.I(WIRE_Data_Cahe_writeData_data[70]), .PAD(PO_Data_Cahe_writeData_data[70]));
PDO02CDG PAD_Data_Cahe_writeData_data71 (.I(WIRE_Data_Cahe_writeData_data[71]), .PAD(PO_Data_Cahe_writeData_data[71]));
PDO02CDG PAD_Data_Cahe_writeData_data72 (.I(WIRE_Data_Cahe_writeData_data[72]), .PAD(PO_Data_Cahe_writeData_data[72]));
PDO02CDG PAD_Data_Cahe_writeData_data73 (.I(WIRE_Data_Cahe_writeData_data[73]), .PAD(PO_Data_Cahe_writeData_data[73]));
PDO02CDG PAD_Data_Cahe_writeData_data74 (.I(WIRE_Data_Cahe_writeData_data[74]), .PAD(PO_Data_Cahe_writeData_data[74]));
PDO02CDG PAD_Data_Cahe_writeData_data75 (.I(WIRE_Data_Cahe_writeData_data[75]), .PAD(PO_Data_Cahe_writeData_data[75]));
PDO02CDG PAD_Data_Cahe_writeData_data76 (.I(WIRE_Data_Cahe_writeData_data[76]), .PAD(PO_Data_Cahe_writeData_data[76]));
PDO02CDG PAD_Data_Cahe_writeData_data77 (.I(WIRE_Data_Cahe_writeData_data[77]), .PAD(PO_Data_Cahe_writeData_data[77]));
PDO02CDG PAD_Data_Cahe_writeData_data78 (.I(WIRE_Data_Cahe_writeData_data[78]), .PAD(PO_Data_Cahe_writeData_data[78]));
PDO02CDG PAD_Data_Cahe_writeData_data79 (.I(WIRE_Data_Cahe_writeData_data[79]), .PAD(PO_Data_Cahe_writeData_data[79]));
PDO02CDG PAD_Data_Cahe_writeData_data80 (.I(WIRE_Data_Cahe_writeData_data[80]), .PAD(PO_Data_Cahe_writeData_data[80]));
PDO02CDG PAD_Data_Cahe_writeData_data81 (.I(WIRE_Data_Cahe_writeData_data[81]), .PAD(PO_Data_Cahe_writeData_data[81]));
PDO02CDG PAD_Data_Cahe_writeData_data82 (.I(WIRE_Data_Cahe_writeData_data[82]), .PAD(PO_Data_Cahe_writeData_data[82]));
PDO02CDG PAD_Data_Cahe_writeData_data83 (.I(WIRE_Data_Cahe_writeData_data[83]), .PAD(PO_Data_Cahe_writeData_data[83]));
PDO02CDG PAD_Data_Cahe_writeData_data84 (.I(WIRE_Data_Cahe_writeData_data[84]), .PAD(PO_Data_Cahe_writeData_data[84]));
PDO02CDG PAD_Data_Cahe_writeData_data85 (.I(WIRE_Data_Cahe_writeData_data[85]), .PAD(PO_Data_Cahe_writeData_data[85]));
PDO02CDG PAD_Data_Cahe_writeData_data86 (.I(WIRE_Data_Cahe_writeData_data[86]), .PAD(PO_Data_Cahe_writeData_data[86]));
PDO02CDG PAD_Data_Cahe_writeData_data87 (.I(WIRE_Data_Cahe_writeData_data[87]), .PAD(PO_Data_Cahe_writeData_data[87]));
PDO02CDG PAD_Data_Cahe_writeData_data88 (.I(WIRE_Data_Cahe_writeData_data[88]), .PAD(PO_Data_Cahe_writeData_data[88]));
PDO02CDG PAD_Data_Cahe_writeData_data89 (.I(WIRE_Data_Cahe_writeData_data[89]), .PAD(PO_Data_Cahe_writeData_data[89]));
PDO02CDG PAD_Data_Cahe_writeData_data90 (.I(WIRE_Data_Cahe_writeData_data[90]), .PAD(PO_Data_Cahe_writeData_data[90]));
PDO02CDG PAD_Data_Cahe_writeData_data91 (.I(WIRE_Data_Cahe_writeData_data[91]), .PAD(PO_Data_Cahe_writeData_data[91]));
PDO02CDG PAD_Data_Cahe_writeData_data92 (.I(WIRE_Data_Cahe_writeData_data[92]), .PAD(PO_Data_Cahe_writeData_data[92]));
PDO02CDG PAD_Data_Cahe_writeData_data93 (.I(WIRE_Data_Cahe_writeData_data[93]), .PAD(PO_Data_Cahe_writeData_data[93]));
PDO02CDG PAD_Data_Cahe_writeData_data94 (.I(WIRE_Data_Cahe_writeData_data[94]), .PAD(PO_Data_Cahe_writeData_data[94]));
PDO02CDG PAD_Data_Cahe_writeData_data95 (.I(WIRE_Data_Cahe_writeData_data[95]), .PAD(PO_Data_Cahe_writeData_data[95]));
PDO02CDG PAD_Data_Cahe_writeData_data96 (.I(WIRE_Data_Cahe_writeData_data[96]), .PAD(PO_Data_Cahe_writeData_data[96]));
PDO02CDG PAD_Data_Cahe_writeData_data97 (.I(WIRE_Data_Cahe_writeData_data[97]), .PAD(PO_Data_Cahe_writeData_data[97]));
PDO02CDG PAD_Data_Cahe_writeData_data98 (.I(WIRE_Data_Cahe_writeData_data[98]), .PAD(PO_Data_Cahe_writeData_data[98]));
PDO02CDG PAD_Data_Cahe_writeData_data99 (.I(WIRE_Data_Cahe_writeData_data[99]), .PAD(PO_Data_Cahe_writeData_data[99]));
PDO02CDG PAD_Data_Cahe_writeData_data100 (.I(WIRE_Data_Cahe_writeData_data[100]), .PAD(PO_Data_Cahe_writeData_data[100]));
PDO02CDG PAD_Data_Cahe_writeData_data101 (.I(WIRE_Data_Cahe_writeData_data[101]), .PAD(PO_Data_Cahe_writeData_data[101]));
PDO02CDG PAD_Data_Cahe_writeData_data102 (.I(WIRE_Data_Cahe_writeData_data[102]), .PAD(PO_Data_Cahe_writeData_data[102]));
PDO02CDG PAD_Data_Cahe_writeData_data103 (.I(WIRE_Data_Cahe_writeData_data[103]), .PAD(PO_Data_Cahe_writeData_data[103]));
PDO02CDG PAD_Data_Cahe_writeData_data104 (.I(WIRE_Data_Cahe_writeData_data[104]), .PAD(PO_Data_Cahe_writeData_data[104]));
PDO02CDG PAD_Data_Cahe_writeData_data105 (.I(WIRE_Data_Cahe_writeData_data[105]), .PAD(PO_Data_Cahe_writeData_data[105]));
PDO02CDG PAD_Data_Cahe_writeData_data106 (.I(WIRE_Data_Cahe_writeData_data[106]), .PAD(PO_Data_Cahe_writeData_data[106]));
PDO02CDG PAD_Data_Cahe_writeData_data107 (.I(WIRE_Data_Cahe_writeData_data[107]), .PAD(PO_Data_Cahe_writeData_data[107]));
PDO02CDG PAD_Data_Cahe_writeData_data108 (.I(WIRE_Data_Cahe_writeData_data[108]), .PAD(PO_Data_Cahe_writeData_data[108]));
PDO02CDG PAD_Data_Cahe_writeData_data109 (.I(WIRE_Data_Cahe_writeData_data[109]), .PAD(PO_Data_Cahe_writeData_data[109]));
PDO02CDG PAD_Data_Cahe_writeData_data110 (.I(WIRE_Data_Cahe_writeData_data[110]), .PAD(PO_Data_Cahe_writeData_data[110]));
PDO02CDG PAD_Data_Cahe_writeData_data111 (.I(WIRE_Data_Cahe_writeData_data[111]), .PAD(PO_Data_Cahe_writeData_data[111]));
PDO02CDG PAD_Data_Cahe_writeData_data112 (.I(WIRE_Data_Cahe_writeData_data[112]), .PAD(PO_Data_Cahe_writeData_data[112]));
PDO02CDG PAD_Data_Cahe_writeData_data113 (.I(WIRE_Data_Cahe_writeData_data[113]), .PAD(PO_Data_Cahe_writeData_data[113]));
PDO02CDG PAD_Data_Cahe_writeData_data114 (.I(WIRE_Data_Cahe_writeData_data[114]), .PAD(PO_Data_Cahe_writeData_data[114]));
PDO02CDG PAD_Data_Cahe_writeData_data115 (.I(WIRE_Data_Cahe_writeData_data[115]), .PAD(PO_Data_Cahe_writeData_data[115]));
PDO02CDG PAD_Data_Cahe_writeData_data116 (.I(WIRE_Data_Cahe_writeData_data[116]), .PAD(PO_Data_Cahe_writeData_data[116]));
PDO02CDG PAD_Data_Cahe_writeData_data117 (.I(WIRE_Data_Cahe_writeData_data[117]), .PAD(PO_Data_Cahe_writeData_data[117]));
PDO02CDG PAD_Data_Cahe_writeData_data118 (.I(WIRE_Data_Cahe_writeData_data[118]), .PAD(PO_Data_Cahe_writeData_data[118]));
PDO02CDG PAD_Data_Cahe_writeData_data119 (.I(WIRE_Data_Cahe_writeData_data[119]), .PAD(PO_Data_Cahe_writeData_data[119]));
PDO02CDG PAD_Data_Cahe_writeData_data120 (.I(WIRE_Data_Cahe_writeData_data[120]), .PAD(PO_Data_Cahe_writeData_data[120]));
PDO02CDG PAD_Data_Cahe_writeData_data121 (.I(WIRE_Data_Cahe_writeData_data[121]), .PAD(PO_Data_Cahe_writeData_data[121]));
PDO02CDG PAD_Data_Cahe_writeData_data122 (.I(WIRE_Data_Cahe_writeData_data[122]), .PAD(PO_Data_Cahe_writeData_data[122]));
PDO02CDG PAD_Data_Cahe_writeData_data123 (.I(WIRE_Data_Cahe_writeData_data[123]), .PAD(PO_Data_Cahe_writeData_data[123]));
PDO02CDG PAD_Data_Cahe_writeData_data124 (.I(WIRE_Data_Cahe_writeData_data[124]), .PAD(PO_Data_Cahe_writeData_data[124]));
PDO02CDG PAD_Data_Cahe_writeData_data125 (.I(WIRE_Data_Cahe_writeData_data[125]), .PAD(PO_Data_Cahe_writeData_data[125]));
PDO02CDG PAD_Data_Cahe_writeData_data126 (.I(WIRE_Data_Cahe_writeData_data[126]), .PAD(PO_Data_Cahe_writeData_data[126]));
PDO02CDG PAD_Data_Cahe_writeData_data127 (.I(WIRE_Data_Cahe_writeData_data[127]), .PAD(PO_Data_Cahe_writeData_data[127]));

PDO02CDG PAD_Data_Cahe_writeData_strb0 (.I(WIRE_Data_Cahe_writeData_strb[0]), .PAD(PO_Data_Cahe_writeData_strb[0]));
PDO02CDG PAD_Data_Cahe_writeData_strb1 (.I(WIRE_Data_Cahe_writeData_strb[1]), .PAD(PO_Data_Cahe_writeData_strb[1]));
PDO02CDG PAD_Data_Cahe_writeData_strb2 (.I(WIRE_Data_Cahe_writeData_strb[2]), .PAD(PO_Data_Cahe_writeData_strb[2]));
PDO02CDG PAD_Data_Cahe_writeData_strb3 (.I(WIRE_Data_Cahe_writeData_strb[3]), .PAD(PO_Data_Cahe_writeData_strb[3]));
PDO02CDG PAD_Data_Cahe_writeData_strb4 (.I(WIRE_Data_Cahe_writeData_strb[4]), .PAD(PO_Data_Cahe_writeData_strb[4]));
PDO02CDG PAD_Data_Cahe_writeData_strb5 (.I(WIRE_Data_Cahe_writeData_strb[5]), .PAD(PO_Data_Cahe_writeData_strb[5]));
PDO02CDG PAD_Data_Cahe_writeData_strb6 (.I(WIRE_Data_Cahe_writeData_strb[6]), .PAD(PO_Data_Cahe_writeData_strb[6]));
PDO02CDG PAD_Data_Cahe_writeData_strb7 (.I(WIRE_Data_Cahe_writeData_strb[7]), .PAD(PO_Data_Cahe_writeData_strb[7]));
PDO02CDG PAD_Data_Cahe_writeData_strb8 (.I(WIRE_Data_Cahe_writeData_strb[8]), .PAD(PO_Data_Cahe_writeData_strb[8]));
PDO02CDG PAD_Data_Cahe_writeData_strb9 (.I(WIRE_Data_Cahe_writeData_strb[9]), .PAD(PO_Data_Cahe_writeData_strb[9]));
PDO02CDG PAD_Data_Cahe_writeData_strb10 (.I(WIRE_Data_Cahe_writeData_strb[10]), .PAD(PO_Data_Cahe_writeData_strb[10]));
PDO02CDG PAD_Data_Cahe_writeData_strb11 (.I(WIRE_Data_Cahe_writeData_strb[11]), .PAD(PO_Data_Cahe_writeData_strb[11]));
PDO02CDG PAD_Data_Cahe_writeData_strb12 (.I(WIRE_Data_Cahe_writeData_strb[12]), .PAD(PO_Data_Cahe_writeData_strb[12]));
PDO02CDG PAD_Data_Cahe_writeData_strb13 (.I(WIRE_Data_Cahe_writeData_strb[13]), .PAD(PO_Data_Cahe_writeData_strb[13]));
PDO02CDG PAD_Data_Cahe_writeData_strb14 (.I(WIRE_Data_Cahe_writeData_strb[14]), .PAD(PO_Data_Cahe_writeData_strb[14]));
PDO02CDG PAD_Data_Cahe_writeData_strb15 (.I(WIRE_Data_Cahe_writeData_strb[15]), .PAD(PO_Data_Cahe_writeData_strb[15]));

PDO02CDG PAD_Data_Cahe_writeData_valid (.I(WIRE_Data_Cahe_writeData_valid), .PAD(PO_Data_Cahe_writeData_valid));
PDO02CDG PAD_Data_Cahe_writeResp_ready (.I(WIRE_Data_Cahe_writeResp_ready), .PAD(PO_Data_Cahe_writeResp_ready));

endmodule


