/*

    AXI Lite 4 Bus
    connecting memory and cache

*/

module AXI_Lite_4_Bus(
    /* IO */
);

// TBD



endmodule